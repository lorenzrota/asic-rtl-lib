../../saci/src/StdRtlPkg.vhd