../../serializer/src/serializer.vhd