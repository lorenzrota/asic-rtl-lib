../../saci/src/saci_master_tb.sv