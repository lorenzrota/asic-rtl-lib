../../12b14benc/src/ssp12b14benc/StdRtlPkg.vhd