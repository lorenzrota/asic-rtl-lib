../../sync/src/sync.vhd