../../saci/src/SaciSlaveRam.vhd