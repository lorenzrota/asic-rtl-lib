* TSMC 13 SACI

.subckt SaciSlave2 rst ack addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] addr[10] addr[11] clk cmd[0] cmd[1] cmd[2] cmd[3] cmd[4] cmd[5] cmd[6] exec rdData[0] rdData[1] rdData[2] rdData[3] rdData[4] rdData[5] rdData[6] rdData[7] rdData[8] rdData[9] rdData[10] rdData[11] rdData[12] rdData[13] rdData[14] rdData[15] rdData[16] rdData[17] rdData[18] rdData[19] rdData[20] rdData[21] rdData[22] rdData[23] rdData[24] rdData[25] rdData[26] rdData[27] rdData[28] rdData[29] rdData[30] rdData[31] readL rstL rstOutL saciCmd saciRsp saciSelL wrData[0] wrData[1] wrData[2] wrData[3] wrData[4] wrData[5] wrData[6] wrData[7] wrData[8] wrData[9] wrData[10] wrData[11] wrData[12] wrData[13] wrData[14] wrData[15] wrData[16] wrData[17] wrData[18] wrData[19] wrData[20] wrData[21] wrData[22] wrData[23] wrData[24] wrData[25] wrData[26] wrData[27] wrData[28] wrData[29] wrData[30] wrData[31]

MU9413/2/1 G_DS CLK U9413/2/2 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-98.32 43.805 -98.19 44.105)
MU9413/2/2 U9413/2/CLK U9413/2/2 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-97.74 43.805 -97.61 44.105)
MU9413/2/3 G_DS CLK U9413/2/3 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-96.56 43.805 -96.43 44.105)
MU9413/2/4 U9413/2/CLK U9413/2/3 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-95.98 43.805 -95.85 44.105)
MU9413/2/5 G_DS U9413/2/CLK U9413/2/4 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-94.8 43.805 -94.67 44.105)
MU9413/2/6 U9413/2/5 U9413/2/4 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-94.22 43.805 -94.09 44.105)
MU9413/2/7 U9413/2/6 U9413/2/ix421/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-93.13 43.805 -93 44.195)
MU9413/2/8 U9413/2/8 U9413/2/5 U9413/2/6 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-92.615 43.805 -92.485 44.195)
MU9413/2/9 U9413/2/9 U9413/2/8 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-91.525 43.805 -91.395 44.105)
MU9413/2/10 U9413/2/10 U9413/2/4 U9413/2/8 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-90.435 43.805 -90.305 44.195)
MU9413/2/11 G_DS U9413/2/CLB U9413/2/10 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-89.815 43.805 -89.685 44.195)
MU9413/2/12 U9413/2/10 U9413/2/9 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-89.195 43.805 -89.065 44.195)
MU9413/2/13 U9413/2/11 U9413/2/9 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-88.105 43.805 -87.975 44.195)
MU9413/2/14 U9413/2/12 U9413/2/4 U9413/2/11 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-87.795 43.805 -87.665 44.195)
MU9413/2/15 U9413/2/13 U9413/2/12 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-86.085 43.805 -85.955 44.105)
MU9413/2/16 U9413/2/14 U9413/2/5 U9413/2/12 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-84.995 43.805 -84.865 44.195)
MU9413/2/17 G_DS U9413/2/CLB U9413/2/14 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-84.415 43.805 -84.285 44.195)
MU9413/2/18 U9413/2/14 U9413/2/13 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-83.835 43.805 -83.705 44.105)
MU9413/2/19 wrData[30] U9413/2/14 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-82.745 43.805 -82.615 44.105)
MU9413/2/20 U9413/2/reg_r_shiftReg_31_/QB U9413/2/13 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-81.655 43.805 -81.525 44.105)
MU9413/2/21 U9413/2/ix421/OUT U9413/2/ix2019/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-80.475 43.805 -80.345 44.065)
MU9413/2/22 G_DS U9413/2/ix2021/OUT U9413/2/ix421/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-79.895 43.805 -79.765 44.065)
MU9413/2/23 U9413/2/20 rdData[30] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-78.715 43.59 -78.585 44.11)
MU9413/2/24 U9413/2/ix2019/OUT wrData[30] U9413/2/20 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-78.135 43.59 -78.005 44.11)
MU9413/2/25 U9413/2/20 U9413/2/ix2019/D U9413/2/ix2019/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-77.555 43.59 -77.425 44.11)
MU9413/2/26 G_DS U9413/2/ix2019/B U9413/2/20 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-76.975 43.59 -76.845 44.11)
MU9413/2/27 U9413/2/ix2021/OUT wrData[29] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-75.795 43.805 -75.665 44.065)
MU9413/2/28 G_DS U9413/2/ix2021/B U9413/2/ix2021/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-75.215 43.805 -75.085 44.065)
MU9413/2/29 U9413/2/29 rdData[29] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-74.035 43.59 -73.905 44.11)
MU9413/2/30 U9413/reg_r_shiftReg_47_\Cross wrData[29] U9413/2/29 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-73.455 43.59 -73.325 44.11)
MU9413/2/31 U9413/2/29 U9413/2/ix2019/D U9413/reg_r_shiftReg_47_\Cross G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-72.875 43.59 -72.745 44.11)
MU9413/2/32 G_DS U9413/2/ix2019/B U9413/2/29 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-72.295 43.59 -72.165 44.11)
MU9413/2/33 G_DS U9413/2/CLK U9413/2/35 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-71.115 43.805 -70.985 44.105)
MU9413/2/34 U9413/2/36 U9413/2/35 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-70.535 43.805 -70.405 44.105)
MU9413/2/35 U9413/2/37 U9413/2/ix397/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-69.445 43.805 -69.315 44.195)
MU9413/2/36 U9413/2/39 U9413/2/36 U9413/2/37 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-68.93 43.805 -68.8 44.195)
MU9413/2/37 U9413/2/40 U9413/2/39 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-67.84 43.805 -67.71 44.105)
MU9413/2/38 U9413/2/41 U9413/2/35 U9413/2/39 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-66.75 43.805 -66.62 44.195)
MU9413/2/39 G_DS U9413/2/CLB U9413/2/41 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-66.13 43.805 -66 44.195)
MU9413/2/40 U9413/2/41 U9413/2/40 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-65.51 43.805 -65.38 44.195)
MU9413/2/41 U9413/2/42 U9413/2/40 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-64.42 43.805 -64.29 44.195)
MU9413/2/42 U9413/2/43 U9413/2/35 U9413/2/42 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-64.11 43.805 -63.98 44.195)
MU9413/2/43 U9413/2/44 U9413/2/43 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-62.4 43.805 -62.27 44.105)
MU9413/2/44 U9413/2/45 U9413/2/36 U9413/2/43 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-61.31 43.805 -61.18 44.195)
MU9413/2/45 G_DS U9413/2/CLB U9413/2/45 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-60.73 43.805 -60.6 44.195)
MU9413/2/46 U9413/2/45 U9413/2/44 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-60.15 43.805 -60.02 44.105)
MU9413/2/47 wrData[28] U9413/2/45 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-59.06 43.805 -58.93 44.105)
MU9413/2/48 U9413/2/reg_r_shiftReg_29_/QB U9413/2/44 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-57.97 43.805 -57.84 44.105)
MU9413/2/49 U9413/2/48 rdData[28] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-56.79 43.59 -56.66 44.11)
MU9413/2/50 U9413/2/ix2031/OUT wrData[28] U9413/2/48 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-56.21 43.59 -56.08 44.11)
MU9413/2/51 U9413/2/48 U9413/2/ix2019/D U9413/2/ix2031/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-55.63 43.59 -55.5 44.11)
MU9413/2/52 G_DS U9413/2/ix2019/B U9413/2/48 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-55.05 43.59 -54.92 44.11)
MU9413/2/53 U9413/2/ix397/OUT U9413/2/ix2031/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-53.87 43.805 -53.74 44.065)
MU9413/2/54 G_DS U9413/2/ix2033/OUT U9413/2/ix397/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-53.29 43.805 -53.16 44.065)
MU9413/2/55 U9413/2/ix2033/OUT wrData[27] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-52.11 43.805 -51.98 44.065)
MU9413/2/56 G_DS U9413/2/ix2021/B U9413/2/ix2033/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-51.53 43.805 -51.4 44.065)
MU9413/2/57 U9413/2/60 rdData[26] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-50.35 43.59 -50.22 44.11)
MU9413/2/58 U9413/2/ix2043/OUT wrData[26] U9413/2/60 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-49.77 43.59 -49.64 44.11)
MU9413/2/59 U9413/2/60 U9413/2/ix2019/D U9413/2/ix2043/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-49.19 43.59 -49.06 44.11)
MU9413/2/60 G_DS U9413/2/ix2019/B U9413/2/60 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-48.61 43.59 -48.48 44.11)
MU9413/2/61 U9413/2/ix373/OUT U9413/2/ix2043/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-47.43 43.805 -47.3 44.065)
MU9413/2/62 G_DS U9413/2/ix2045/OUT U9413/2/ix373/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-46.85 43.805 -46.72 44.065)
MU9413/2/63 U9413/2/ix2045/OUT wrData[25] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-45.67 43.805 -45.54 44.065)
MU9413/2/64 G_DS U9413/2/ix2045/B U9413/2/ix2045/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-45.09 43.805 -44.96 44.065)
MU9413/2/65 U9413/2/ix2051/OUT wrData[24] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-43.91 43.805 -43.78 44.065)
MU9413/2/66 G_DS U9413/2/ix2045/B U9413/2/ix2051/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-43.33 43.805 -43.2 44.065)
MU9413/2/67 U9413/2/ix361/OUT U9413/2/ix2049/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-42.15 43.805 -42.02 44.065)
MU9413/2/68 G_DS U9413/2/ix2051/OUT U9413/2/ix361/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-41.57 43.805 -41.44 44.065)
MU9413/2/69 U9413/2/78 rdData[25] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-40.39 43.59 -40.26 44.11)
MU9413/2/70 U9413/2/ix2049/OUT wrData[25] U9413/2/78 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-39.81 43.59 -39.68 44.11)
MU9413/2/71 U9413/2/78 U9413/2/ix2019/D U9413/2/ix2049/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-39.23 43.59 -39.1 44.11)
MU9413/2/72 G_DS U9413/2/ix2019/B U9413/2/78 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-38.65 43.59 -38.52 44.11)
MU9413/2/73 G_DS U9413/2/CLK U9413/2/84 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-37.47 43.805 -37.34 44.105)
MU9413/2/74 U9413/2/85 U9413/2/84 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-36.89 43.805 -36.76 44.105)
MU9413/2/75 U9413/2/86 U9413/2/ix361/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-35.8 43.805 -35.67 44.195)
MU9413/2/76 U9413/2/88 U9413/2/85 U9413/2/86 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-35.285 43.805 -35.155 44.195)
MU9413/2/77 U9413/2/89 U9413/2/88 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-34.195 43.805 -34.065 44.105)
MU9413/2/78 U9413/2/90 U9413/2/84 U9413/2/88 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-33.105 43.805 -32.975 44.195)
MU9413/2/79 G_DS U9413/2/CLB U9413/2/90 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-32.485 43.805 -32.355 44.195)
MU9413/2/80 U9413/2/90 U9413/2/89 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-31.865 43.805 -31.735 44.195)
MU9413/2/81 U9413/2/91 U9413/2/89 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-30.775 43.805 -30.645 44.195)
MU9413/2/82 U9413/2/92 U9413/2/84 U9413/2/91 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-30.465 43.805 -30.335 44.195)
MU9413/2/83 U9413/2/93 U9413/2/92 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-28.755 43.805 -28.625 44.105)
MU9413/2/84 U9413/2/94 U9413/2/85 U9413/2/92 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-27.665 43.805 -27.535 44.195)
MU9413/2/85 G_DS U9413/2/CLB U9413/2/94 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-27.085 43.805 -26.955 44.195)
MU9413/2/86 U9413/2/94 U9413/2/93 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-26.505 43.805 -26.375 44.105)
MU9413/2/87 wrData[25] U9413/2/94 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-25.415 43.805 -25.285 44.105)
MU9413/2/88 U9413/2/reg_r_shiftReg_26_/QB U9413/2/93 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-24.325 43.805 -24.195 44.105)
MU9413/2/89 U9413/2/97 rdData[23] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-23.145 43.59 -23.015 44.11)
MU9413/2/90 U9413/2/ix2061/OUT wrData[23] U9413/2/97 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-22.565 43.59 -22.435 44.11)
MU9413/2/91 U9413/2/97 U9413/2/ix2019/D U9413/2/ix2061/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-21.985 43.59 -21.855 44.11)
MU9413/2/92 G_DS U9413/2/ix2019/B U9413/2/97 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-21.405 43.59 -21.275 44.11)
MU9413/2/93 G_DS U9413/2/CLK U9413/2/103 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-20.225 43.805 -20.095 44.105)
MU9413/2/94 U9413/2/104 U9413/2/103 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-19.645 43.805 -19.515 44.105)
MU9413/2/95 U9413/2/105 U9413/2/ix325/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-18.555 43.805 -18.425 44.195)
MU9413/2/96 U9413/2/107 U9413/2/104 U9413/2/105 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-18.04 43.805 -17.91 44.195)
MU9413/2/97 U9413/2/108 U9413/2/107 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-16.95 43.805 -16.82 44.105)
MU9413/2/98 U9413/2/109 U9413/2/103 U9413/2/107 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-15.86 43.805 -15.73 44.195)
MU9413/2/99 G_DS U9413/2/CLB U9413/2/109 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-15.24 43.805 -15.11 44.195)
MU9413/2/100 U9413/2/109 U9413/2/108 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-14.62 43.805 -14.49 44.195)
MU9413/2/101 U9413/2/110 U9413/2/108 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-13.53 43.805 -13.4 44.195)
MU9413/2/102 U9413/2/111 U9413/2/103 U9413/2/110 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-13.22 43.805 -13.09 44.195)
MU9413/2/103 U9413/2/112 U9413/2/111 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-11.51 43.805 -11.38 44.105)
MU9413/2/104 U9413/2/113 U9413/2/104 U9413/2/111 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-10.42 43.805 -10.29 44.195)
MU9413/2/105 G_DS U9413/2/CLB U9413/2/113 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-9.84 43.805 -9.71 44.195)
MU9413/2/106 U9413/2/113 U9413/2/112 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-9.26 43.805 -9.13 44.105)
MU9413/2/107 wrData[22] U9413/2/113 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-8.17 43.805 -8.04 44.105)
MU9413/2/108 U9413/2/reg_r_shiftReg_23_/QB U9413/2/112 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-7.08 43.805 -6.95 44.105)
MU9413/2/109 U9413/2/116 rdData[22] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-5.9 43.59 -5.77 44.11)
MU9413/2/110 U9413/2/ix2067/OUT wrData[22] U9413/2/116 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-5.32 43.59 -5.19 44.11)
MU9413/2/111 U9413/2/116 U9413/2/ix2067/D U9413/2/ix2067/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-4.74 43.59 -4.61 44.11)
MU9413/2/112 G_DS U9413/2/ix2067/B U9413/2/116 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-4.16 43.59 -4.03 44.11)
MU9413/2/113 U9413/2/ix325/OUT U9413/2/ix2067/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-2.98 43.805 -2.85 44.065)
MU9413/2/114 G_DS U9413/2/ix2069/OUT U9413/2/ix325/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-2.4 43.805 -2.27 44.065)
MU9413/2/115 U9413/2/ix2069/OUT wrData[21] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-1.22 43.805 -1.09 44.065)
MU9413/2/116 G_DS U9413/2/ix2045/B U9413/2/ix2069/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-0.64 43.805 -0.51 44.065)
MU9413/2/117 U9413/2/128 rdData[20] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(0.54 43.59 0.67 44.11)
MU9413/2/118 U9413/2/ix2079/OUT wrData[20] U9413/2/128 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(1.12 43.59 1.25 44.11)
MU9413/2/119 U9413/2/128 U9413/2/ix2067/D U9413/2/ix2079/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(1.7 43.59 1.83 44.11)
MU9413/2/120 G_DS U9413/2/ix2067/B U9413/2/128 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(2.28 43.59 2.41 44.11)
MU9413/2/121 U9413/2/134 rdData[19] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(3.46 43.59 3.59 44.11)
MU9413/2/122 U9413/2/ix2085/OUT wrData[19] U9413/2/134 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(4.04 43.59 4.17 44.11)
MU9413/2/123 U9413/2/134 U9413/2/ix2067/D U9413/2/ix2085/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(4.62 43.59 4.75 44.11)
MU9413/2/124 G_DS U9413/2/ix2067/B U9413/2/134 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(5.2 43.59 5.33 44.11)
MU9413/2/125 U9413/2/ix289/OUT U9413/2/ix2085/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(6.38 43.805 6.51 44.065)
MU9413/2/126 G_DS U9413/2/ix2087/OUT U9413/2/ix289/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(6.96 43.805 7.09 44.065)
MU9413/2/127 U9413/2/ix2087/OUT wrData[18] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(8.14 43.805 8.27 44.065)
MU9413/2/128 G_DS U9413/2/ix2045/B U9413/2/ix2087/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(8.72 43.805 8.85 44.065)
MU9413/2/129 U9413/2/146 rdData[18] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(9.9 43.59 10.03 44.11)
MU9413/2/130 U9413/2/ix2091/OUT wrData[18] U9413/2/146 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(10.48 43.59 10.61 44.11)
MU9413/2/131 U9413/2/146 U9413/2/ix2067/D U9413/2/ix2091/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(11.06 43.59 11.19 44.11)
MU9413/2/132 G_DS U9413/2/ix2067/B U9413/2/146 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(11.64 43.59 11.77 44.11)
MU9413/2/133 U9413/2/ix277/OUT U9413/2/ix2091/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(12.82 43.805 12.95 44.065)
MU9413/2/134 G_DS U9413/2/ix2093/OUT U9413/2/ix277/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(13.4 43.805 13.53 44.065)
MU9413/2/135 U9413/2/ix2093/OUT wrData[17] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(14.58 43.805 14.71 44.065)
MU9413/2/136 G_DS U9413/2/ix2093/B U9413/2/ix2093/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(15.16 43.805 15.29 44.065)
MU9413/2/137 G_DS U9413/2/CLK U9413/2/158 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(16.34 43.805 16.47 44.105)
MU9413/2/138 U9413/2/159 U9413/2/158 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(16.92 43.805 17.05 44.105)
MU9413/2/139 U9413/2/160 U9413/2/ix277/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(18.01 43.805 18.14 44.195)
MU9413/2/140 U9413/2/162 U9413/2/159 U9413/2/160 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(18.525 43.805 18.655 44.195)
MU9413/2/141 U9413/2/163 U9413/2/162 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(19.615 43.805 19.745 44.105)
MU9413/2/142 U9413/2/164 U9413/2/158 U9413/2/162 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(20.705 43.805 20.835 44.195)
MU9413/2/143 G_DS U9413/2/CLB U9413/2/164 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(21.325 43.805 21.455 44.195)
MU9413/2/144 U9413/2/164 U9413/2/163 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(21.945 43.805 22.075 44.195)
MU9413/2/145 U9413/2/165 U9413/2/163 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(23.035 43.805 23.165 44.195)
MU9413/2/146 U9413/2/166 U9413/2/158 U9413/2/165 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(23.345 43.805 23.475 44.195)
MU9413/2/147 U9413/2/167 U9413/2/166 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(25.055 43.805 25.185 44.105)
MU9413/2/148 U9413/2/168 U9413/2/159 U9413/2/166 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(26.145 43.805 26.275 44.195)
MU9413/2/149 G_DS U9413/2/CLB U9413/2/168 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(26.725 43.805 26.855 44.195)
MU9413/2/150 U9413/2/168 U9413/2/167 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(27.305 43.805 27.435 44.105)
MU9413/2/151 wrData[18] U9413/2/168 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(28.395 43.805 28.525 44.105)
MU9413/2/152 U9413/2/reg_r_shiftReg_19_/QB U9413/2/167 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(29.485 43.805 29.615 44.105)
MU9413/2/153 U9413/2/ix2105/OUT wrData[15] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(30.665 43.805 30.795 44.065)
MU9413/2/154 G_DS U9413/2/ix2093/B U9413/2/ix2105/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(31.245 43.805 31.375 44.065)
MU9413/2/155 U9413/2/174 rdData[15] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(32.425 43.59 32.555 44.11)
MU9413/2/156 U9413/2/ix2109/OUT wrData[15] U9413/2/174 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(33.005 43.59 33.135 44.11)
MU9413/2/157 U9413/2/174 U9413/2/ix2067/D U9413/2/ix2109/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(33.585 43.59 33.715 44.11)
MU9413/2/158 G_DS U9413/2/ix2067/B U9413/2/174 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(34.165 43.59 34.295 44.11)
MU9413/2/159 U9413/2/ix241/OUT U9413/2/ix2109/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(35.345 43.805 35.475 44.065)
MU9413/2/160 G_DS U9413/2/ix2111/OUT U9413/2/ix241/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(35.925 43.805 36.055 44.065)
MU9413/2/161 U9413/2/ix2111/OUT wrData[14] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(37.105 43.805 37.235 44.065)
MU9413/2/162 G_DS U9413/2/ix2093/B U9413/2/ix2111/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(37.685 43.805 37.815 44.065)
MU9413/2/163 G_DS U9413/2/CLK U9413/2/186 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(38.865 43.805 38.995 44.105)
MU9413/2/164 U9413/2/187 U9413/2/186 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(39.445 43.805 39.575 44.105)
MU9413/2/165 U9413/2/188 U9413/2/ix241/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(40.535 43.805 40.665 44.195)
MU9413/2/166 U9413/2/190 U9413/2/187 U9413/2/188 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(41.05 43.805 41.18 44.195)
MU9413/2/167 U9413/2/191 U9413/2/190 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(42.14 43.805 42.27 44.105)
MU9413/2/168 U9413/2/192 U9413/2/186 U9413/2/190 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(43.23 43.805 43.36 44.195)
MU9413/2/169 G_DS U9413/2/CLB U9413/2/192 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(43.85 43.805 43.98 44.195)
MU9413/2/170 U9413/2/192 U9413/2/191 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(44.47 43.805 44.6 44.195)
MU9413/2/171 U9413/2/193 U9413/2/191 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(45.56 43.805 45.69 44.195)
MU9413/2/172 U9413/2/194 U9413/2/186 U9413/2/193 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(45.87 43.805 46 44.195)
MU9413/2/173 U9413/2/195 U9413/2/194 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(47.58 43.805 47.71 44.105)
MU9413/2/174 U9413/2/196 U9413/2/187 U9413/2/194 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(48.67 43.805 48.8 44.195)
MU9413/2/175 G_DS U9413/2/CLB U9413/2/196 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(49.25 43.805 49.38 44.195)
MU9413/2/176 U9413/2/196 U9413/2/195 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(49.83 43.805 49.96 44.105)
MU9413/2/177 wrData[15] U9413/2/196 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(50.92 43.805 51.05 44.105)
MU9413/2/178 U9413/2/reg_r_shiftReg_16_/QB U9413/2/195 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(52.01 43.805 52.14 44.105)
MU9413/2/179 U9413/2/199 rdData[13] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(53.19 43.59 53.32 44.11)
MU9413/2/180 U9413/2/ix2121/OUT wrData[13] U9413/2/199 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(53.77 43.59 53.9 44.11)
MU9413/2/181 U9413/2/199 U9413/2/ix2121/D U9413/2/ix2121/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(54.35 43.59 54.48 44.11)
MU9413/2/182 G_DS U9413/2/ix2121/B U9413/2/199 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(54.93 43.59 55.06 44.11)
MU9413/2/183 U9413/2/205 rdData[12] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(56.11 43.59 56.24 44.11)
MU9413/2/184 U9413/2/ix2127/OUT wrData[12] U9413/2/205 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(56.69 43.59 56.82 44.11)
MU9413/2/185 U9413/2/205 U9413/2/ix2121/D U9413/2/ix2127/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(57.27 43.59 57.4 44.11)
MU9413/2/186 G_DS U9413/2/ix2121/B U9413/2/205 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(57.85 43.59 57.98 44.11)
MU9413/2/187 U9413/2/211 rdData[11] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(59.03 43.59 59.16 44.11)
MU9413/2/188 U9413/2/ix2133/OUT wrData[11] U9413/2/211 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(59.61 43.59 59.74 44.11)
MU9413/2/189 U9413/2/211 U9413/2/ix2121/D U9413/2/ix2133/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(60.19 43.59 60.32 44.11)
MU9413/2/190 G_DS U9413/2/ix2121/B U9413/2/211 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(60.77 43.59 60.9 44.11)
MU9413/2/191 U9413/2/ix181/B wrData[9] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(61.95 43.805 62.08 44.065)
MU9413/2/192 G_DS U9413/2/ix2093/B U9413/2/ix181/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(62.53 43.805 62.66 44.065)
MU9413/2/193 U9413/2/ix181/OUT U9413/2/ix181/A G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(63.71 43.805 63.84 44.065)
MU9413/2/194 G_DS U9413/2/ix181/B U9413/2/ix181/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(64.29 43.805 64.42 44.065)
MU9413/2/195 U9413/2/223 rdData[10] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(65.47 43.59 65.6 44.11)
MU9413/2/196 U9413/2/ix181/A wrData[10] U9413/2/223 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(66.05 43.59 66.18 44.11)
MU9413/2/197 U9413/2/223 U9413/2/ix2121/D U9413/2/ix181/A G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(66.63 43.59 66.76 44.11)
MU9413/2/198 G_DS U9413/2/ix2121/B U9413/2/223 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(67.21 43.59 67.34 44.11)
MU9413/2/199 U9413/2/ix169/B wrData[8] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(68.39 43.805 68.52 44.065)
MU9413/2/200 G_DS U9413/2/ix2147/B U9413/2/ix169/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(68.97 43.805 69.1 44.065)
MU9413/2/201 U9413/2/ix169/OUT U9413/2/ix169/A G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(70.15 43.805 70.28 44.065)
MU9413/2/202 G_DS U9413/2/ix169/B U9413/2/ix169/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(70.73 43.805 70.86 44.065)
MU9413/2/203 U9413/2/235 rdData[9] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(71.91 43.59 72.04 44.11)
MU9413/2/204 U9413/2/ix169/A wrData[9] U9413/2/235 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(72.49 43.59 72.62 44.11)
MU9413/2/205 U9413/2/235 U9413/2/ix2121/D U9413/2/ix169/A G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(73.07 43.59 73.2 44.11)
MU9413/2/206 G_DS U9413/2/ix2121/B U9413/2/235 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(73.65 43.59 73.78 44.11)
MU9413/2/207 G_DS U9413/2/CLK U9413/2/241 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(74.83 43.805 74.96 44.105)
MU9413/2/208 U9413/2/242 U9413/2/241 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(75.41 43.805 75.54 44.105)
MU9413/2/209 U9413/2/243 U9413/2/ix169/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(76.5 43.805 76.63 44.195)
MU9413/2/210 U9413/2/245 U9413/2/242 U9413/2/243 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(77.015 43.805 77.145 44.195)
MU9413/2/211 U9413/2/246 U9413/2/245 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(78.105 43.805 78.235 44.105)
MU9413/2/212 U9413/2/247 U9413/2/241 U9413/2/245 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(79.195 43.805 79.325 44.195)
MU9413/2/213 G_DS U9413/2/CLB U9413/2/247 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(79.815 43.805 79.945 44.195)
MU9413/2/214 U9413/2/247 U9413/2/246 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(80.435 43.805 80.565 44.195)
MU9413/2/215 U9413/2/248 U9413/2/246 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(81.525 43.805 81.655 44.195)
MU9413/2/216 U9413/2/249 U9413/2/241 U9413/2/248 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(81.835 43.805 81.965 44.195)
MU9413/2/217 U9413/2/250 U9413/2/249 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(83.545 43.805 83.675 44.105)
MU9413/2/218 U9413/2/251 U9413/2/242 U9413/2/249 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(84.635 43.805 84.765 44.195)
MU9413/2/219 G_DS U9413/2/CLB U9413/2/251 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(85.215 43.805 85.345 44.195)
MU9413/2/220 U9413/2/251 U9413/2/250 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(85.795 43.805 85.925 44.105)
MU9413/2/221 wrData[9] U9413/2/251 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(86.885 43.805 87.015 44.105)
MU9413/2/222 U9413/2/reg_r_shiftReg_10_/QB U9413/2/250 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(87.975 43.805 88.105 44.105)
MU9413/2/223 U9413/2/254 rdData[5] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(89.155 43.59 89.285 44.11)
MU9413/2/224 U9413/2/ix121/A wrData[5] U9413/2/254 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(89.735 43.59 89.865 44.11)
MU9413/2/225 U9413/2/254 U9413/2/ix2121/D U9413/2/ix121/A G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(90.315 43.59 90.445 44.11)
MU9413/2/226 G_DS U9413/2/ix2121/B U9413/2/254 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(90.895 43.59 91.025 44.11)
MU9413/2/227 U9413/2/ix121/OUT U9413/2/ix121/A G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(92.075 43.805 92.205 44.065)
MU9413/2/228 G_DS U9413/2/ix121/B U9413/2/ix121/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(92.655 43.805 92.785 44.065)
MU9413/2/229 U9413/2/ix121/B wrData[4] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(93.835 43.805 93.965 44.065)
MU9413/2/230 G_DS U9413/2/ix2147/B U9413/2/ix121/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(94.415 43.805 94.545 44.065)
MU9413/2/231 G_DS U9413/2/CLK U9413/2/266 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(95.595 43.805 95.725 44.105)
MU9413/2/232 U9413/2/267 U9413/2/266 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(96.175 43.805 96.305 44.105)
MU9413/2/233 U9413/2/268 U9413/2/ix121/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(97.265 43.805 97.395 44.195)
MU9413/2/234 U9413/2/270 U9413/2/267 U9413/2/268 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(97.78 43.805 97.91 44.195)
MU9413/2/235 U9413/2/271 U9413/2/270 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(98.87 43.805 99 44.105)
MU9413/2/236 U9413/2/272 U9413/2/266 U9413/2/270 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(99.96 43.805 100.09 44.195)
MU9413/2/237 G_DS U9413/2/CLB U9413/2/272 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(100.58 43.805 100.71 44.195)
MU9413/2/238 U9413/2/272 U9413/2/271 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(101.2 43.805 101.33 44.195)
MU9413/2/239 U9413/2/273 U9413/2/271 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(102.29 43.805 102.42 44.195)
MU9413/2/240 U9413/2/274 U9413/2/266 U9413/2/273 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(102.6 43.805 102.73 44.195)
MU9413/2/241 U9413/2/275 U9413/2/274 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(104.31 43.805 104.44 44.105)
MU9413/2/242 U9413/2/276 U9413/2/267 U9413/2/274 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(105.4 43.805 105.53 44.195)
MU9413/2/243 G_DS U9413/2/CLB U9413/2/276 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(105.98 43.805 106.11 44.195)
MU9413/2/244 U9413/2/276 U9413/2/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(106.56 43.805 106.69 44.105)
MU9413/2/245 wrData[5] U9413/2/276 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(107.65 43.805 107.78 44.105)
MU9413/2/246 U9413/2/reg_r_shiftReg_6_/QB U9413/2/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(108.74 43.805 108.87 44.105)
MU9413/2/247 U9413/2/279 rdData[4] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(109.92 43.59 110.05 44.11)
MU9413/2/248 U9413/2/ix2175/OUT wrData[4] U9413/2/279 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(110.5 43.59 110.63 44.11)
MU9413/2/249 U9413/2/279 U9413/D U9413/2/ix2175/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(111.08 43.59 111.21 44.11)
MU9413/2/250 G_DS U9413/2/ix1948/B U9413/2/279 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(111.66 43.59 111.79 44.11)
MU9413/2/251 U9413/2/ix2189/OUT wrData[1] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(112.84 43.805 112.97 44.065)
MU9413/2/252 G_DS U9413/2/ix2147/B U9413/2/ix2189/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(113.42 43.805 113.55 44.065)
MU9413/2/253 U9413/2/ix61/OUT U9413/2/ix1948/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(114.6 43.805 114.73 44.065)
MU9413/2/254 G_DS U9413/reg_r_shiftReg_21_\Cross U9413/2/ix61/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(115.18 43.805 115.31 44.065)
MU9413/2/255 G_DS U9413/2/CLK U9413/2/291 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(116.36 43.805 116.49 44.105)
MU9413/2/256 U9413/2/292 U9413/2/291 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(116.94 43.805 117.07 44.105)
MU9413/2/257 U9413/2/293 U9413/2/ix61/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(118.03 43.805 118.16 44.195)
MU9413/2/258 U9413/2/295 U9413/2/292 U9413/2/293 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(118.545 43.805 118.675 44.195)
MU9413/2/259 U9413/2/296 U9413/2/295 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(119.635 43.805 119.765 44.105)
MU9413/2/260 U9413/2/297 U9413/2/291 U9413/2/295 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(120.725 43.805 120.855 44.195)
MU9413/2/261 G_DS U9413/2/CLB U9413/2/297 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(121.345 43.805 121.475 44.195)
MU9413/2/262 U9413/2/297 U9413/2/296 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(121.965 43.805 122.095 44.195)
MU9413/2/263 U9413/2/298 U9413/2/296 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(123.055 43.805 123.185 44.195)
MU9413/2/264 U9413/2/299 U9413/2/291 U9413/2/298 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(123.365 43.805 123.495 44.195)
MU9413/2/265 U9413/2/300 U9413/2/299 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(125.075 43.805 125.205 44.105)
MU9413/2/266 U9413/2/301 U9413/2/292 U9413/2/299 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(126.165 43.805 126.295 44.195)
MU9413/2/267 G_DS U9413/2/CLB U9413/2/301 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(126.745 43.805 126.875 44.195)
MU9413/2/268 U9413/2/301 U9413/2/300 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(127.325 43.805 127.455 44.105)
MU9413/2/269 wrData[0] U9413/2/301 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(128.415 43.805 128.545 44.105)
MU9413/2/270 U9413/2/reg_r_shiftReg_1_/QB U9413/2/300 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(129.505 43.805 129.635 44.105)
MU9413/2/271 U9413/2/304 rdData[0] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(130.685 43.59 130.815 44.11)
MU9413/2/272 U9413/2/ix1948/OUT wrData[0] U9413/2/304 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(131.265 43.59 131.395 44.11)
MU9413/2/273 U9413/2/304 U9413/D U9413/2/ix1948/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(131.845 43.59 131.975 44.11)
MU9413/2/274 G_DS U9413/2/ix1948/B U9413/2/304 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(132.425 43.59 132.555 44.11)
MU9413/2/275 U9413/2/310 rdData[1] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(133.605 43.59 133.735 44.11)
MU9413/2/276 U9413/2/ix2193/OUT wrData[1] U9413/2/310 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(134.185 43.59 134.315 44.11)
MU9413/2/277 U9413/2/310 U9413/D U9413/2/ix2193/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(134.765 43.59 134.895 44.11)
MU9413/2/278 G_DS U9413/2/ix1948/B U9413/2/310 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(135.345 43.59 135.475 44.11)
MU9413/2/279 U9413/2/ix2195/OUT wrData[0] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(136.525 43.805 136.655 44.065)
MU9413/2/280 G_DS U9413/2/ix2147/B U9413/2/ix2195/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(137.105 43.805 137.235 44.065)
MU9413/2/281 U9413/DATA U9413/2/ix2193/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(138.285 43.805 138.415 44.065)
MU9413/2/282 G_DS U9413/2/ix2195/OUT U9413/DATA G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(138.865 43.805 138.995 44.065)
MU9413/2/283 G_DS U9413/2/CLK U9413/2/320 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(140.045 43.805 140.175 44.105)
MU9413/2/284 U9413/2/321 U9413/2/320 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(140.625 43.805 140.755 44.105)
MU9413/2/285 U9413/2/322 U9413/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(141.715 43.805 141.845 44.195)
MU9413/2/286 U9413/2/323 U9413/2/321 U9413/2/322 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(142.23 43.805 142.36 44.195)
MU9413/2/287 U9413/2/324 U9413/2/323 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(143.32 43.805 143.45 44.105)
MU9413/2/288 U9413/2/325 U9413/2/320 U9413/2/323 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(144.41 43.805 144.54 44.195)
MU9413/2/289 G_DS U9413/2/CLB U9413/2/325 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(145.03 43.805 145.16 44.195)
MU9413/2/290 U9413/2/325 U9413/2/324 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(145.65 43.805 145.78 44.195)
MU9413/2/291 U9413/2/326 U9413/2/324 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(146.74 43.805 146.87 44.195)
MU9413/2/292 U9413/2/327 U9413/2/320 U9413/2/326 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(147.05 43.805 147.18 44.195)
MU9413/2/293 U9413/2/328 U9413/2/327 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(148.76 43.805 148.89 44.105)
MU9413/2/294 U9413/2/329 U9413/2/321 U9413/2/327 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(149.85 43.805 149.98 44.195)
MU9413/2/295 G_DS U9413/2/CLB U9413/2/329 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(150.43 43.805 150.56 44.195)
MU9413/2/296 U9413/2/329 U9413/2/328 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(151.01 43.805 151.14 44.105)
MU9413/2/297 wrData[1] U9413/2/329 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(152.1 43.805 152.23 44.105)
MU9413/2/298 U9413/2/reg_r_shiftReg_2_/QB U9413/2/328 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(153.19 43.805 153.32 44.105)
MU9413/2/299 U9413/2/331 U9413/OUT G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(154.37 43.59 154.5 44.11)
MU9413/2/300 RST saciSelL U9413/2/331 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(154.95 43.59 155.08 44.11)
MU9413/2/301 U9413/OUT rstL G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(156.13 43.805 156.26 44.105)
MU9413/2/302 G_DS RST U9413/2/334 G_DS pch sa=-3.65e-007 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(157.31 43.805 157.44 44.105)
MU9413/2/303 U9413/2/CLB U9413/2/334 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(157.89 43.805 158.02 44.105)
MU9413/2/304 G_DS RST U9413/2/335 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(159.07 43.805 159.2 44.105)
MU9413/2/305 U9413/2/CLB U9413/2/335 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(159.65 43.805 159.78 44.105)
MU9413/2/right_51/1 G_DG RST U9413/2/334 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(157.31 42.075 157.44 42.225)
MU9413/2/right_51/2 U9413/2/CLB U9413/2/334 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(157.89 42.075 158.02 42.225)
MU9413/2/right_50/1 G_DG RST U9413/2/335 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(159.07 42.075 159.2 42.225)
MU9413/2/right_50/2 U9413/2/CLB U9413/2/335 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(159.65 42.075 159.78 42.225)
MU9413/2/left_51/1 G_DG CLK U9413/2/2 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-98.32 42.075 -98.19 42.225)
MU9413/2/left_51/2 U9413/2/CLK U9413/2/2 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-97.74 42.075 -97.61 42.225)
MU9413/2/left_50/1 G_DG CLK U9413/2/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-96.56 42.075 -96.43 42.225)
MU9413/2/left_50/2 U9413/2/CLK U9413/2/3 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-95.98 42.075 -95.85 42.225)
MU9413/2/ix2259/1 U9413/OUT rstL G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(156.13 42.075 156.26 42.225)
MU9413/2/ix499/1 RST U9413/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(154.37 42.075 154.5 42.225)
MU9413/2/ix499/2 G_DG saciSelL RST G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(154.95 42.075 155.08 42.225)
MU9413/2/reg_r_shiftReg_2_/1 G_DG U9413/2/CLK U9413/2/320 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(140.045 42.075 140.175 42.225)
MU9413/2/reg_r_shiftReg_2_/2 U9413/2/321 U9413/2/320 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(140.625 42.075 140.755 42.225)
MU9413/2/reg_r_shiftReg_2_/3 U9413/2/reg_r_shiftReg_2_/4 U9413/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(141.715 42.075 141.845 42.225)
MU9413/2/reg_r_shiftReg_2_/4 U9413/2/323 U9413/2/320 U9413/2/reg_r_shiftReg_2_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(142.23 42.075 142.36 42.225)
MU9413/2/reg_r_shiftReg_2_/5 U9413/2/324 U9413/2/323 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(143.32 42.075 143.45 42.225)
MU9413/2/reg_r_shiftReg_2_/6 U9413/2/reg_r_shiftReg_2_/7 U9413/2/CLB U9413/2/323 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(144.69 42.075 144.82 42.225)
MU9413/2/reg_r_shiftReg_2_/7 U9413/2/reg_r_shiftReg_2_/8 U9413/2/324 U9413/2/reg_r_shiftReg_2_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(145.17 42.075 145.3 42.225)
MU9413/2/reg_r_shiftReg_2_/8 G_DG U9413/2/321 U9413/2/reg_r_shiftReg_2_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(145.65 42.075 145.78 42.225)
MU9413/2/reg_r_shiftReg_2_/9 U9413/2/reg_r_shiftReg_2_/9 U9413/2/324 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(146.74 42.075 146.87 42.225)
MU9413/2/reg_r_shiftReg_2_/10 U9413/2/reg_r_shiftReg_2_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_2_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(147.25 42.075 147.38 42.225)
MU9413/2/reg_r_shiftReg_2_/11 U9413/2/327 U9413/2/321 U9413/2/reg_r_shiftReg_2_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(147.67 42.075 147.8 42.225)
MU9413/2/reg_r_shiftReg_2_/12 U9413/2/328 U9413/2/327 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(148.76 42.075 148.89 42.225)
MU9413/2/reg_r_shiftReg_2_/13 U9413/2/329 U9413/2/320 U9413/2/327 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(150.12 42.075 150.25 42.225)
MU9413/2/reg_r_shiftReg_2_/14 U9413/2/reg_r_shiftReg_2_/14 U9413/2/CLB U9413/2/329 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(150.7 42.075 150.83 42.225)
MU9413/2/reg_r_shiftReg_2_/15 G_DG U9413/2/328 U9413/2/reg_r_shiftReg_2_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(151.01 42.075 151.14 42.225)
MU9413/2/reg_r_shiftReg_2_/16 wrData[1] U9413/2/329 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(152.1 42.075 152.23 42.225)
MU9413/2/reg_r_shiftReg_2_/17 U9413/2/reg_r_shiftReg_2_/QB U9413/2/328 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(153.19 42.075 153.32 42.225)
MU9413/2/ix73/1 U9413/2/ix73/1 U9413/2/ix2193/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(138.285 42.075 138.415 42.225)
MU9413/2/ix73/2 U9413/DATA U9413/2/ix2195/OUT U9413/2/ix73/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(138.865 42.075 138.995 42.225)
MU9413/2/ix2195/1 U9413/2/ix2195/1 wrData[0] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(136.525 42.075 136.655 42.225)
MU9413/2/ix2195/2 U9413/2/ix2195/OUT U9413/2/ix2147/B U9413/2/ix2195/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(137.105 42.075 137.235 42.225)
MU9413/2/ix2193/1 U9413/2/ix2193/1 rdData[1] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(133.605 42.075 133.735 42.225)
MU9413/2/ix2193/2 U9413/2/ix2193/OUT U9413/2/ix1948/B U9413/2/ix2193/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(134.185 42.075 134.315 42.225)
MU9413/2/ix2193/3 U9413/2/ix2193/3 wrData[1] U9413/2/ix2193/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(134.765 42.075 134.895 42.225)
MU9413/2/ix2193/4 G_DG U9413/D U9413/2/ix2193/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(135.345 42.075 135.475 42.225)
MU9413/2/ix1948/1 U9413/2/ix1948/1 rdData[0] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(130.685 42.075 130.815 42.225)
MU9413/2/ix1948/2 U9413/2/ix1948/OUT U9413/2/ix1948/B U9413/2/ix1948/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(131.265 42.075 131.395 42.225)
MU9413/2/ix1948/3 U9413/2/ix1948/3 wrData[0] U9413/2/ix1948/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(131.845 42.075 131.975 42.225)
MU9413/2/ix1948/4 G_DG U9413/D U9413/2/ix1948/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(132.425 42.075 132.555 42.225)
MU9413/2/reg_r_shiftReg_1_/1 G_DG U9413/2/CLK U9413/2/291 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(116.36 42.075 116.49 42.225)
MU9413/2/reg_r_shiftReg_1_/2 U9413/2/292 U9413/2/291 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(116.94 42.075 117.07 42.225)
MU9413/2/reg_r_shiftReg_1_/3 U9413/2/reg_r_shiftReg_1_/4 U9413/2/ix61/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(118.03 42.075 118.16 42.225)
MU9413/2/reg_r_shiftReg_1_/4 U9413/2/295 U9413/2/291 U9413/2/reg_r_shiftReg_1_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(118.545 42.075 118.675 42.225)
MU9413/2/reg_r_shiftReg_1_/5 U9413/2/296 U9413/2/295 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(119.635 42.075 119.765 42.225)
MU9413/2/reg_r_shiftReg_1_/6 U9413/2/reg_r_shiftReg_1_/7 U9413/2/CLB U9413/2/295 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(121.005 42.075 121.135 42.225)
MU9413/2/reg_r_shiftReg_1_/7 U9413/2/reg_r_shiftReg_1_/8 U9413/2/296 U9413/2/reg_r_shiftReg_1_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(121.485 42.075 121.615 42.225)
MU9413/2/reg_r_shiftReg_1_/8 G_DG U9413/2/292 U9413/2/reg_r_shiftReg_1_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(121.965 42.075 122.095 42.225)
MU9413/2/reg_r_shiftReg_1_/9 U9413/2/reg_r_shiftReg_1_/9 U9413/2/296 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(123.055 42.075 123.185 42.225)
MU9413/2/reg_r_shiftReg_1_/10 U9413/2/reg_r_shiftReg_1_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_1_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(123.565 42.075 123.695 42.225)
MU9413/2/reg_r_shiftReg_1_/11 U9413/2/299 U9413/2/292 U9413/2/reg_r_shiftReg_1_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(123.985 42.075 124.115 42.225)
MU9413/2/reg_r_shiftReg_1_/12 U9413/2/300 U9413/2/299 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(125.075 42.075 125.205 42.225)
MU9413/2/reg_r_shiftReg_1_/13 U9413/2/301 U9413/2/291 U9413/2/299 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(126.435 42.075 126.565 42.225)
MU9413/2/reg_r_shiftReg_1_/14 U9413/2/reg_r_shiftReg_1_/14 U9413/2/CLB U9413/2/301 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(127.015 42.075 127.145 42.225)
MU9413/2/reg_r_shiftReg_1_/15 G_DG U9413/2/300 U9413/2/reg_r_shiftReg_1_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(127.325 42.075 127.455 42.225)
MU9413/2/reg_r_shiftReg_1_/16 wrData[0] U9413/2/301 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(128.415 42.075 128.545 42.225)
MU9413/2/reg_r_shiftReg_1_/17 U9413/2/reg_r_shiftReg_1_/QB U9413/2/300 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(129.505 42.075 129.635 42.225)
MU9413/2/ix61/1 U9413/2/ix61/1 U9413/2/ix1948/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(114.6 42.075 114.73 42.225)
MU9413/2/ix61/2 U9413/2/ix61/OUT U9413/reg_r_shiftReg_21_\Cross U9413/2/ix61/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(115.18 42.075 115.31 42.225)
MU9413/2/ix2189/1 U9413/2/ix2189/1 wrData[1] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(112.84 42.075 112.97 42.225)
MU9413/2/ix2189/2 U9413/2/ix2189/OUT U9413/2/ix2147/B U9413/2/ix2189/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(113.42 42.075 113.55 42.225)
MU9413/2/ix2175/1 U9413/2/ix2175/1 rdData[4] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(109.92 42.075 110.05 42.225)
MU9413/2/ix2175/2 U9413/2/ix2175/OUT U9413/2/ix1948/B U9413/2/ix2175/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(110.5 42.075 110.63 42.225)
MU9413/2/ix2175/3 U9413/2/ix2175/3 wrData[4] U9413/2/ix2175/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(111.08 42.075 111.21 42.225)
MU9413/2/ix2175/4 G_DG U9413/D U9413/2/ix2175/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(111.66 42.075 111.79 42.225)
MU9413/2/reg_r_shiftReg_6_/1 G_DG U9413/2/CLK U9413/2/266 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(95.595 42.075 95.725 42.225)
MU9413/2/reg_r_shiftReg_6_/2 U9413/2/267 U9413/2/266 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(96.175 42.075 96.305 42.225)
MU9413/2/reg_r_shiftReg_6_/3 U9413/2/reg_r_shiftReg_6_/4 U9413/2/ix121/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(97.265 42.075 97.395 42.225)
MU9413/2/reg_r_shiftReg_6_/4 U9413/2/270 U9413/2/266 U9413/2/reg_r_shiftReg_6_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(97.78 42.075 97.91 42.225)
MU9413/2/reg_r_shiftReg_6_/5 U9413/2/271 U9413/2/270 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(98.87 42.075 99 42.225)
MU9413/2/reg_r_shiftReg_6_/6 U9413/2/reg_r_shiftReg_6_/7 U9413/2/CLB U9413/2/270 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(100.24 42.075 100.37 42.225)
MU9413/2/reg_r_shiftReg_6_/7 U9413/2/reg_r_shiftReg_6_/8 U9413/2/271 U9413/2/reg_r_shiftReg_6_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(100.72 42.075 100.85 42.225)
MU9413/2/reg_r_shiftReg_6_/8 G_DG U9413/2/267 U9413/2/reg_r_shiftReg_6_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(101.2 42.075 101.33 42.225)
MU9413/2/reg_r_shiftReg_6_/9 U9413/2/reg_r_shiftReg_6_/9 U9413/2/271 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(102.29 42.075 102.42 42.225)
MU9413/2/reg_r_shiftReg_6_/10 U9413/2/reg_r_shiftReg_6_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_6_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(102.8 42.075 102.93 42.225)
MU9413/2/reg_r_shiftReg_6_/11 U9413/2/274 U9413/2/267 U9413/2/reg_r_shiftReg_6_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(103.22 42.075 103.35 42.225)
MU9413/2/reg_r_shiftReg_6_/12 U9413/2/275 U9413/2/274 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(104.31 42.075 104.44 42.225)
MU9413/2/reg_r_shiftReg_6_/13 U9413/2/276 U9413/2/266 U9413/2/274 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(105.67 42.075 105.8 42.225)
MU9413/2/reg_r_shiftReg_6_/14 U9413/2/reg_r_shiftReg_6_/14 U9413/2/CLB U9413/2/276 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(106.25 42.075 106.38 42.225)
MU9413/2/reg_r_shiftReg_6_/15 G_DG U9413/2/275 U9413/2/reg_r_shiftReg_6_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(106.56 42.075 106.69 42.225)
MU9413/2/reg_r_shiftReg_6_/16 wrData[5] U9413/2/276 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(107.65 42.075 107.78 42.225)
MU9413/2/reg_r_shiftReg_6_/17 U9413/2/reg_r_shiftReg_6_/QB U9413/2/275 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(108.74 42.075 108.87 42.225)
MU9413/2/ix2171/1 U9413/2/ix2171/1 wrData[4] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(93.835 42.075 93.965 42.225)
MU9413/2/ix2171/2 U9413/2/ix121/B U9413/2/ix2147/B U9413/2/ix2171/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(94.415 42.075 94.545 42.225)
MU9413/2/ix121/1 U9413/2/ix121/1 U9413/2/ix121/A G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(92.075 42.075 92.205 42.225)
MU9413/2/ix121/2 U9413/2/ix121/OUT U9413/2/ix121/B U9413/2/ix121/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(92.655 42.075 92.785 42.225)
MU9413/2/ix2169/1 U9413/2/ix2169/1 rdData[5] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(89.155 42.075 89.285 42.225)
MU9413/2/ix2169/2 U9413/2/ix121/A U9413/2/ix2121/B U9413/2/ix2169/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(89.735 42.075 89.865 42.225)
MU9413/2/ix2169/3 U9413/2/ix2169/3 wrData[5] U9413/2/ix121/A G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(90.315 42.075 90.445 42.225)
MU9413/2/ix2169/4 G_DG U9413/2/ix2121/D U9413/2/ix2169/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(90.895 42.075 91.025 42.225)
MU9413/2/reg_r_shiftReg_10_/1 G_DG U9413/2/CLK U9413/2/241 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(74.83 42.075 74.96 42.225)
MU9413/2/reg_r_shiftReg_10_/2 U9413/2/242 U9413/2/241 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(75.41 42.075 75.54 42.225)
MU9413/2/reg_r_shiftReg_10_/3 U9413/2/reg_r_shiftReg_10_/4 U9413/2/ix169/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(76.5 42.075 76.63 42.225)
MU9413/2/reg_r_shiftReg_10_/4 U9413/2/245 U9413/2/241 U9413/2/reg_r_shiftReg_10_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(77.015 42.075 77.145 42.225)
MU9413/2/reg_r_shiftReg_10_/5 U9413/2/246 U9413/2/245 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(78.105 42.075 78.235 42.225)
MU9413/2/reg_r_shiftReg_10_/6 U9413/2/reg_r_shiftReg_10_/7 U9413/2/CLB U9413/2/245 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(79.475 42.075 79.605 42.225)
MU9413/2/reg_r_shiftReg_10_/7 U9413/2/reg_r_shiftReg_10_/8 U9413/2/246 U9413/2/reg_r_shiftReg_10_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(79.955 42.075 80.085 42.225)
MU9413/2/reg_r_shiftReg_10_/8 G_DG U9413/2/242 U9413/2/reg_r_shiftReg_10_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(80.435 42.075 80.565 42.225)
MU9413/2/reg_r_shiftReg_10_/9 U9413/2/reg_r_shiftReg_10_/9 U9413/2/246 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(81.525 42.075 81.655 42.225)
MU9413/2/reg_r_shiftReg_10_/10 U9413/2/reg_r_shiftReg_10_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_10_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(82.035 42.075 82.165 42.225)
MU9413/2/reg_r_shiftReg_10_/11 U9413/2/249 U9413/2/242 U9413/2/reg_r_shiftReg_10_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(82.455 42.075 82.585 42.225)
MU9413/2/reg_r_shiftReg_10_/12 U9413/2/250 U9413/2/249 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(83.545 42.075 83.675 42.225)
MU9413/2/reg_r_shiftReg_10_/13 U9413/2/251 U9413/2/241 U9413/2/249 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(84.905 42.075 85.035 42.225)
MU9413/2/reg_r_shiftReg_10_/14 U9413/2/reg_r_shiftReg_10_/14 U9413/2/CLB U9413/2/251 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(85.485 42.075 85.615 42.225)
MU9413/2/reg_r_shiftReg_10_/15 G_DG U9413/2/250 U9413/2/reg_r_shiftReg_10_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(85.795 42.075 85.925 42.225)
MU9413/2/reg_r_shiftReg_10_/16 wrData[9] U9413/2/251 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(86.885 42.075 87.015 42.225)
MU9413/2/reg_r_shiftReg_10_/17 U9413/2/reg_r_shiftReg_10_/QB U9413/2/250 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(87.975 42.075 88.105 42.225)
MU9413/2/ix2145/1 U9413/2/ix2145/1 rdData[9] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(71.91 42.075 72.04 42.225)
MU9413/2/ix2145/2 U9413/2/ix169/A U9413/2/ix2121/B U9413/2/ix2145/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(72.49 42.075 72.62 42.225)
MU9413/2/ix2145/3 U9413/2/ix2145/3 wrData[9] U9413/2/ix169/A G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(73.07 42.075 73.2 42.225)
MU9413/2/ix2145/4 G_DG U9413/2/ix2121/D U9413/2/ix2145/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(73.65 42.075 73.78 42.225)
MU9413/2/ix169/1 U9413/2/ix169/1 U9413/2/ix169/A G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(70.15 42.075 70.28 42.225)
MU9413/2/ix169/2 U9413/2/ix169/OUT U9413/2/ix169/B U9413/2/ix169/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(70.73 42.075 70.86 42.225)
MU9413/2/ix2147/1 U9413/2/ix2147/1 wrData[8] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(68.39 42.075 68.52 42.225)
MU9413/2/ix2147/2 U9413/2/ix169/B U9413/2/ix2147/B U9413/2/ix2147/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(68.97 42.075 69.1 42.225)
MU9413/2/ix2139/1 U9413/2/ix2139/1 rdData[10] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(65.47 42.075 65.6 42.225)
MU9413/2/ix2139/2 U9413/2/ix181/A U9413/2/ix2121/B U9413/2/ix2139/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(66.05 42.075 66.18 42.225)
MU9413/2/ix2139/3 U9413/2/ix2139/3 wrData[10] U9413/2/ix181/A G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(66.63 42.075 66.76 42.225)
MU9413/2/ix2139/4 G_DG U9413/2/ix2121/D U9413/2/ix2139/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(67.21 42.075 67.34 42.225)
MU9413/2/ix181/1 U9413/2/ix181/1 U9413/2/ix181/A G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(63.71 42.075 63.84 42.225)
MU9413/2/ix181/2 U9413/2/ix181/OUT U9413/2/ix181/B U9413/2/ix181/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(64.29 42.075 64.42 42.225)
MU9413/2/ix2141/1 U9413/2/ix2141/1 wrData[9] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(61.95 42.075 62.08 42.225)
MU9413/2/ix2141/2 U9413/2/ix181/B U9413/2/ix2093/B U9413/2/ix2141/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(62.53 42.075 62.66 42.225)
MU9413/2/ix2133/1 U9413/2/ix2133/1 rdData[11] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(59.03 42.075 59.16 42.225)
MU9413/2/ix2133/2 U9413/2/ix2133/OUT U9413/2/ix2121/B U9413/2/ix2133/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(59.61 42.075 59.74 42.225)
MU9413/2/ix2133/3 U9413/2/ix2133/3 wrData[11] U9413/2/ix2133/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(60.19 42.075 60.32 42.225)
MU9413/2/ix2133/4 G_DG U9413/2/ix2121/D U9413/2/ix2133/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(60.77 42.075 60.9 42.225)
MU9413/2/ix2127/1 U9413/2/ix2127/1 rdData[12] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(56.11 42.075 56.24 42.225)
MU9413/2/ix2127/2 U9413/2/ix2127/OUT U9413/2/ix2121/B U9413/2/ix2127/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(56.69 42.075 56.82 42.225)
MU9413/2/ix2127/3 U9413/2/ix2127/3 wrData[12] U9413/2/ix2127/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(57.27 42.075 57.4 42.225)
MU9413/2/ix2127/4 G_DG U9413/2/ix2121/D U9413/2/ix2127/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(57.85 42.075 57.98 42.225)
MU9413/2/ix2121/1 U9413/2/ix2121/1 rdData[13] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(53.19 42.075 53.32 42.225)
MU9413/2/ix2121/2 U9413/2/ix2121/OUT U9413/2/ix2121/B U9413/2/ix2121/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(53.77 42.075 53.9 42.225)
MU9413/2/ix2121/3 U9413/2/ix2121/3 wrData[13] U9413/2/ix2121/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(54.35 42.075 54.48 42.225)
MU9413/2/ix2121/4 G_DG U9413/2/ix2121/D U9413/2/ix2121/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(54.93 42.075 55.06 42.225)
MU9413/2/reg_r_shiftReg_16_/1 G_DG U9413/2/CLK U9413/2/186 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(38.865 42.075 38.995 42.225)
MU9413/2/reg_r_shiftReg_16_/2 U9413/2/187 U9413/2/186 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(39.445 42.075 39.575 42.225)
MU9413/2/reg_r_shiftReg_16_/3 U9413/2/reg_r_shiftReg_16_/4 U9413/2/ix241/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(40.535 42.075 40.665 42.225)
MU9413/2/reg_r_shiftReg_16_/4 U9413/2/190 U9413/2/186 U9413/2/reg_r_shiftReg_16_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(41.05 42.075 41.18 42.225)
MU9413/2/reg_r_shiftReg_16_/5 U9413/2/191 U9413/2/190 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(42.14 42.075 42.27 42.225)
MU9413/2/reg_r_shiftReg_16_/6 U9413/2/reg_r_shiftReg_16_/7 U9413/2/CLB U9413/2/190 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(43.51 42.075 43.64 42.225)
MU9413/2/reg_r_shiftReg_16_/7 U9413/2/reg_r_shiftReg_16_/8 U9413/2/191 U9413/2/reg_r_shiftReg_16_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(43.99 42.075 44.12 42.225)
MU9413/2/reg_r_shiftReg_16_/8 G_DG U9413/2/187 U9413/2/reg_r_shiftReg_16_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(44.47 42.075 44.6 42.225)
MU9413/2/reg_r_shiftReg_16_/9 U9413/2/reg_r_shiftReg_16_/9 U9413/2/191 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(45.56 42.075 45.69 42.225)
MU9413/2/reg_r_shiftReg_16_/10 U9413/2/reg_r_shiftReg_16_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_16_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(46.07 42.075 46.2 42.225)
MU9413/2/reg_r_shiftReg_16_/11 U9413/2/194 U9413/2/187 U9413/2/reg_r_shiftReg_16_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(46.49 42.075 46.62 42.225)
MU9413/2/reg_r_shiftReg_16_/12 U9413/2/195 U9413/2/194 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(47.58 42.075 47.71 42.225)
MU9413/2/reg_r_shiftReg_16_/13 U9413/2/196 U9413/2/186 U9413/2/194 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(48.94 42.075 49.07 42.225)
MU9413/2/reg_r_shiftReg_16_/14 U9413/2/reg_r_shiftReg_16_/14 U9413/2/CLB U9413/2/196 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(49.52 42.075 49.65 42.225)
MU9413/2/reg_r_shiftReg_16_/15 G_DG U9413/2/195 U9413/2/reg_r_shiftReg_16_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(49.83 42.075 49.96 42.225)
MU9413/2/reg_r_shiftReg_16_/16 wrData[15] U9413/2/196 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(50.92 42.075 51.05 42.225)
MU9413/2/reg_r_shiftReg_16_/17 U9413/2/reg_r_shiftReg_16_/QB U9413/2/195 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(52.01 42.075 52.14 42.225)
MU9413/2/ix2111/1 U9413/2/ix2111/1 wrData[14] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(37.105 42.075 37.235 42.225)
MU9413/2/ix2111/2 U9413/2/ix2111/OUT U9413/2/ix2093/B U9413/2/ix2111/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(37.685 42.075 37.815 42.225)
MU9413/2/ix241/1 U9413/2/ix241/1 U9413/2/ix2109/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(35.345 42.075 35.475 42.225)
MU9413/2/ix241/2 U9413/2/ix241/OUT U9413/2/ix2111/OUT U9413/2/ix241/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(35.925 42.075 36.055 42.225)
MU9413/2/ix2109/1 U9413/2/ix2109/1 rdData[15] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(32.425 42.075 32.555 42.225)
MU9413/2/ix2109/2 U9413/2/ix2109/OUT U9413/2/ix2067/B U9413/2/ix2109/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(33.005 42.075 33.135 42.225)
MU9413/2/ix2109/3 U9413/2/ix2109/3 wrData[15] U9413/2/ix2109/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(33.585 42.075 33.715 42.225)
MU9413/2/ix2109/4 G_DG U9413/2/ix2067/D U9413/2/ix2109/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(34.165 42.075 34.295 42.225)
MU9413/2/ix2105/1 U9413/2/ix2105/1 wrData[15] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(30.665 42.075 30.795 42.225)
MU9413/2/ix2105/2 U9413/2/ix2105/OUT U9413/2/ix2093/B U9413/2/ix2105/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(31.245 42.075 31.375 42.225)
MU9413/2/reg_r_shiftReg_19_/1 G_DG U9413/2/CLK U9413/2/158 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(16.34 42.075 16.47 42.225)
MU9413/2/reg_r_shiftReg_19_/2 U9413/2/159 U9413/2/158 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(16.92 42.075 17.05 42.225)
MU9413/2/reg_r_shiftReg_19_/3 U9413/2/reg_r_shiftReg_19_/4 U9413/2/ix277/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(18.01 42.075 18.14 42.225)
MU9413/2/reg_r_shiftReg_19_/4 U9413/2/162 U9413/2/158 U9413/2/reg_r_shiftReg_19_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(18.525 42.075 18.655 42.225)
MU9413/2/reg_r_shiftReg_19_/5 U9413/2/163 U9413/2/162 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(19.615 42.075 19.745 42.225)
MU9413/2/reg_r_shiftReg_19_/6 U9413/2/reg_r_shiftReg_19_/7 U9413/2/CLB U9413/2/162 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(20.985 42.075 21.115 42.225)
MU9413/2/reg_r_shiftReg_19_/7 U9413/2/reg_r_shiftReg_19_/8 U9413/2/163 U9413/2/reg_r_shiftReg_19_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(21.465 42.075 21.595 42.225)
MU9413/2/reg_r_shiftReg_19_/8 G_DG U9413/2/159 U9413/2/reg_r_shiftReg_19_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(21.945 42.075 22.075 42.225)
MU9413/2/reg_r_shiftReg_19_/9 U9413/2/reg_r_shiftReg_19_/9 U9413/2/163 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(23.035 42.075 23.165 42.225)
MU9413/2/reg_r_shiftReg_19_/10 U9413/2/reg_r_shiftReg_19_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_19_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(23.545 42.075 23.675 42.225)
MU9413/2/reg_r_shiftReg_19_/11 U9413/2/166 U9413/2/159 U9413/2/reg_r_shiftReg_19_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(23.965 42.075 24.095 42.225)
MU9413/2/reg_r_shiftReg_19_/12 U9413/2/167 U9413/2/166 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(25.055 42.075 25.185 42.225)
MU9413/2/reg_r_shiftReg_19_/13 U9413/2/168 U9413/2/158 U9413/2/166 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(26.415 42.075 26.545 42.225)
MU9413/2/reg_r_shiftReg_19_/14 U9413/2/reg_r_shiftReg_19_/14 U9413/2/CLB U9413/2/168 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(26.995 42.075 27.125 42.225)
MU9413/2/reg_r_shiftReg_19_/15 G_DG U9413/2/167 U9413/2/reg_r_shiftReg_19_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(27.305 42.075 27.435 42.225)
MU9413/2/reg_r_shiftReg_19_/16 wrData[18] U9413/2/168 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(28.395 42.075 28.525 42.225)
MU9413/2/reg_r_shiftReg_19_/17 U9413/2/reg_r_shiftReg_19_/QB U9413/2/167 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(29.485 42.075 29.615 42.225)
MU9413/2/ix2093/1 U9413/2/ix2093/1 wrData[17] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(14.58 42.075 14.71 42.225)
MU9413/2/ix2093/2 U9413/2/ix2093/OUT U9413/2/ix2093/B U9413/2/ix2093/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(15.16 42.075 15.29 42.225)
MU9413/2/ix277/1 U9413/2/ix277/1 U9413/2/ix2091/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(12.82 42.075 12.95 42.225)
MU9413/2/ix277/2 U9413/2/ix277/OUT U9413/2/ix2093/OUT U9413/2/ix277/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(13.4 42.075 13.53 42.225)
MU9413/2/ix2091/1 U9413/2/ix2091/1 rdData[18] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(9.9 42.075 10.03 42.225)
MU9413/2/ix2091/2 U9413/2/ix2091/OUT U9413/2/ix2067/B U9413/2/ix2091/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(10.48 42.075 10.61 42.225)
MU9413/2/ix2091/3 U9413/2/ix2091/3 wrData[18] U9413/2/ix2091/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(11.06 42.075 11.19 42.225)
MU9413/2/ix2091/4 G_DG U9413/2/ix2067/D U9413/2/ix2091/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(11.64 42.075 11.77 42.225)
MU9413/2/ix2087/1 U9413/2/ix2087/1 wrData[18] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(8.14 42.075 8.27 42.225)
MU9413/2/ix2087/2 U9413/2/ix2087/OUT U9413/2/ix2045/B U9413/2/ix2087/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(8.72 42.075 8.85 42.225)
MU9413/2/ix289/1 U9413/2/ix289/1 U9413/2/ix2085/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(6.38 42.075 6.51 42.225)
MU9413/2/ix289/2 U9413/2/ix289/OUT U9413/2/ix2087/OUT U9413/2/ix289/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(6.96 42.075 7.09 42.225)
MU9413/2/ix2085/1 U9413/2/ix2085/1 rdData[19] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(3.46 42.075 3.59 42.225)
MU9413/2/ix2085/2 U9413/2/ix2085/OUT U9413/2/ix2067/B U9413/2/ix2085/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(4.04 42.075 4.17 42.225)
MU9413/2/ix2085/3 U9413/2/ix2085/3 wrData[19] U9413/2/ix2085/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(4.62 42.075 4.75 42.225)
MU9413/2/ix2085/4 G_DG U9413/2/ix2067/D U9413/2/ix2085/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(5.2 42.075 5.33 42.225)
MU9413/2/ix2079/1 U9413/2/ix2079/1 rdData[20] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(0.54 42.075 0.67 42.225)
MU9413/2/ix2079/2 U9413/2/ix2079/OUT U9413/2/ix2067/B U9413/2/ix2079/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(1.12 42.075 1.25 42.225)
MU9413/2/ix2079/3 U9413/2/ix2079/3 wrData[20] U9413/2/ix2079/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(1.7 42.075 1.83 42.225)
MU9413/2/ix2079/4 G_DG U9413/2/ix2067/D U9413/2/ix2079/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(2.28 42.075 2.41 42.225)
MU9413/2/ix2069/1 U9413/2/ix2069/1 wrData[21] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-1.22 42.075 -1.09 42.225)
MU9413/2/ix2069/2 U9413/2/ix2069/OUT U9413/2/ix2045/B U9413/2/ix2069/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-0.64 42.075 -0.51 42.225)
MU9413/2/ix325/1 U9413/2/ix325/1 U9413/2/ix2067/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-2.98 42.075 -2.85 42.225)
MU9413/2/ix325/2 U9413/2/ix325/OUT U9413/2/ix2069/OUT U9413/2/ix325/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-2.4 42.075 -2.27 42.225)
MU9413/2/ix2067/1 U9413/2/ix2067/1 rdData[22] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-5.9 42.075 -5.77 42.225)
MU9413/2/ix2067/2 U9413/2/ix2067/OUT U9413/2/ix2067/B U9413/2/ix2067/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-5.32 42.075 -5.19 42.225)
MU9413/2/ix2067/3 U9413/2/ix2067/3 wrData[22] U9413/2/ix2067/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-4.74 42.075 -4.61 42.225)
MU9413/2/ix2067/4 G_DG U9413/2/ix2067/D U9413/2/ix2067/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-4.16 42.075 -4.03 42.225)
MU9413/2/reg_r_shiftReg_23_/1 G_DG U9413/2/CLK U9413/2/103 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-20.225 42.075 -20.095 42.225)
MU9413/2/reg_r_shiftReg_23_/2 U9413/2/104 U9413/2/103 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-19.645 42.075 -19.515 42.225)
MU9413/2/reg_r_shiftReg_23_/3 U9413/2/reg_r_shiftReg_23_/4 U9413/2/ix325/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-18.555 42.075 -18.425 42.225)
MU9413/2/reg_r_shiftReg_23_/4 U9413/2/107 U9413/2/103 U9413/2/reg_r_shiftReg_23_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-18.04 42.075 -17.91 42.225)
MU9413/2/reg_r_shiftReg_23_/5 U9413/2/108 U9413/2/107 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-16.95 42.075 -16.82 42.225)
MU9413/2/reg_r_shiftReg_23_/6 U9413/2/reg_r_shiftReg_23_/7 U9413/2/CLB U9413/2/107 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-15.58 42.075 -15.45 42.225)
MU9413/2/reg_r_shiftReg_23_/7 U9413/2/reg_r_shiftReg_23_/8 U9413/2/108 U9413/2/reg_r_shiftReg_23_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-15.1 42.075 -14.97 42.225)
MU9413/2/reg_r_shiftReg_23_/8 G_DG U9413/2/104 U9413/2/reg_r_shiftReg_23_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-14.62 42.075 -14.49 42.225)
MU9413/2/reg_r_shiftReg_23_/9 U9413/2/reg_r_shiftReg_23_/9 U9413/2/108 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-13.53 42.075 -13.4 42.225)
MU9413/2/reg_r_shiftReg_23_/10 U9413/2/reg_r_shiftReg_23_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_23_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-13.02 42.075 -12.89 42.225)
MU9413/2/reg_r_shiftReg_23_/11 U9413/2/111 U9413/2/104 U9413/2/reg_r_shiftReg_23_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-12.6 42.075 -12.47 42.225)
MU9413/2/reg_r_shiftReg_23_/12 U9413/2/112 U9413/2/111 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-11.51 42.075 -11.38 42.225)
MU9413/2/reg_r_shiftReg_23_/13 U9413/2/113 U9413/2/103 U9413/2/111 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-10.15 42.075 -10.02 42.225)
MU9413/2/reg_r_shiftReg_23_/14 U9413/2/reg_r_shiftReg_23_/14 U9413/2/CLB U9413/2/113 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-9.57 42.075 -9.44 42.225)
MU9413/2/reg_r_shiftReg_23_/15 G_DG U9413/2/112 U9413/2/reg_r_shiftReg_23_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-9.26 42.075 -9.13 42.225)
MU9413/2/reg_r_shiftReg_23_/16 wrData[22] U9413/2/113 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-8.17 42.075 -8.04 42.225)
MU9413/2/reg_r_shiftReg_23_/17 U9413/2/reg_r_shiftReg_23_/QB U9413/2/112 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-7.08 42.075 -6.95 42.225)
MU9413/2/ix2061/1 U9413/2/ix2061/1 rdData[23] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-23.145 42.075 -23.015 42.225)
MU9413/2/ix2061/2 U9413/2/ix2061/OUT U9413/2/ix2019/B U9413/2/ix2061/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-22.565 42.075 -22.435 42.225)
MU9413/2/ix2061/3 U9413/2/ix2061/3 wrData[23] U9413/2/ix2061/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-21.985 42.075 -21.855 42.225)
MU9413/2/ix2061/4 G_DG U9413/2/ix2019/D U9413/2/ix2061/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-21.405 42.075 -21.275 42.225)
MU9413/2/reg_r_shiftReg_26_/1 G_DG U9413/2/CLK U9413/2/84 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-37.47 42.075 -37.34 42.225)
MU9413/2/reg_r_shiftReg_26_/2 U9413/2/85 U9413/2/84 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-36.89 42.075 -36.76 42.225)
MU9413/2/reg_r_shiftReg_26_/3 U9413/2/reg_r_shiftReg_26_/4 U9413/2/ix361/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-35.8 42.075 -35.67 42.225)
MU9413/2/reg_r_shiftReg_26_/4 U9413/2/88 U9413/2/84 U9413/2/reg_r_shiftReg_26_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-35.285 42.075 -35.155 42.225)
MU9413/2/reg_r_shiftReg_26_/5 U9413/2/89 U9413/2/88 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-34.195 42.075 -34.065 42.225)
MU9413/2/reg_r_shiftReg_26_/6 U9413/2/reg_r_shiftReg_26_/7 U9413/2/CLB U9413/2/88 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-32.825 42.075 -32.695 42.225)
MU9413/2/reg_r_shiftReg_26_/7 U9413/2/reg_r_shiftReg_26_/8 U9413/2/89 U9413/2/reg_r_shiftReg_26_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-32.345 42.075 -32.215 42.225)
MU9413/2/reg_r_shiftReg_26_/8 G_DG U9413/2/85 U9413/2/reg_r_shiftReg_26_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-31.865 42.075 -31.735 42.225)
MU9413/2/reg_r_shiftReg_26_/9 U9413/2/reg_r_shiftReg_26_/9 U9413/2/89 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-30.775 42.075 -30.645 42.225)
MU9413/2/reg_r_shiftReg_26_/10 U9413/2/reg_r_shiftReg_26_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_26_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-30.265 42.075 -30.135 42.225)
MU9413/2/reg_r_shiftReg_26_/11 U9413/2/92 U9413/2/85 U9413/2/reg_r_shiftReg_26_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-29.845 42.075 -29.715 42.225)
MU9413/2/reg_r_shiftReg_26_/12 U9413/2/93 U9413/2/92 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-28.755 42.075 -28.625 42.225)
MU9413/2/reg_r_shiftReg_26_/13 U9413/2/94 U9413/2/84 U9413/2/92 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-27.395 42.075 -27.265 42.225)
MU9413/2/reg_r_shiftReg_26_/14 U9413/2/reg_r_shiftReg_26_/14 U9413/2/CLB U9413/2/94 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-26.815 42.075 -26.685 42.225)
MU9413/2/reg_r_shiftReg_26_/15 G_DG U9413/2/93 U9413/2/reg_r_shiftReg_26_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-26.505 42.075 -26.375 42.225)
MU9413/2/reg_r_shiftReg_26_/16 wrData[25] U9413/2/94 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-25.415 42.075 -25.285 42.225)
MU9413/2/reg_r_shiftReg_26_/17 U9413/2/reg_r_shiftReg_26_/QB U9413/2/93 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-24.325 42.075 -24.195 42.225)
MU9413/2/ix2049/1 U9413/2/ix2049/1 rdData[25] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-40.39 42.075 -40.26 42.225)
MU9413/2/ix2049/2 U9413/2/ix2049/OUT U9413/2/ix2019/B U9413/2/ix2049/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-39.81 42.075 -39.68 42.225)
MU9413/2/ix2049/3 U9413/2/ix2049/3 wrData[25] U9413/2/ix2049/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-39.23 42.075 -39.1 42.225)
MU9413/2/ix2049/4 G_DG U9413/2/ix2019/D U9413/2/ix2049/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-38.65 42.075 -38.52 42.225)
MU9413/2/ix361/1 U9413/2/ix361/1 U9413/2/ix2049/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-42.15 42.075 -42.02 42.225)
MU9413/2/ix361/2 U9413/2/ix361/OUT U9413/2/ix2051/OUT U9413/2/ix361/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-41.57 42.075 -41.44 42.225)
MU9413/2/ix2051/1 U9413/2/ix2051/1 wrData[24] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-43.91 42.075 -43.78 42.225)
MU9413/2/ix2051/2 U9413/2/ix2051/OUT U9413/2/ix2045/B U9413/2/ix2051/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-43.33 42.075 -43.2 42.225)
MU9413/2/ix2045/1 U9413/2/ix2045/1 wrData[25] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-45.67 42.075 -45.54 42.225)
MU9413/2/ix2045/2 U9413/2/ix2045/OUT U9413/2/ix2045/B U9413/2/ix2045/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-45.09 42.075 -44.96 42.225)
MU9413/2/ix373/1 U9413/2/ix373/1 U9413/2/ix2043/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-47.43 42.075 -47.3 42.225)
MU9413/2/ix373/2 U9413/2/ix373/OUT U9413/2/ix2045/OUT U9413/2/ix373/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-46.85 42.075 -46.72 42.225)
MU9413/2/ix2043/1 U9413/2/ix2043/1 rdData[26] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-50.35 42.075 -50.22 42.225)
MU9413/2/ix2043/2 U9413/2/ix2043/OUT U9413/2/ix2019/B U9413/2/ix2043/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-49.77 42.075 -49.64 42.225)
MU9413/2/ix2043/3 U9413/2/ix2043/3 wrData[26] U9413/2/ix2043/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-49.19 42.075 -49.06 42.225)
MU9413/2/ix2043/4 G_DG U9413/2/ix2019/D U9413/2/ix2043/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-48.61 42.075 -48.48 42.225)
MU9413/2/ix2033/1 U9413/2/ix2033/1 wrData[27] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-52.11 42.075 -51.98 42.225)
MU9413/2/ix2033/2 U9413/2/ix2033/OUT U9413/2/ix2021/B U9413/2/ix2033/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-51.53 42.075 -51.4 42.225)
MU9413/2/ix397/1 U9413/2/ix397/1 U9413/2/ix2031/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-53.87 42.075 -53.74 42.225)
MU9413/2/ix397/2 U9413/2/ix397/OUT U9413/2/ix2033/OUT U9413/2/ix397/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-53.29 42.075 -53.16 42.225)
MU9413/2/ix2031/1 U9413/2/ix2031/1 rdData[28] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-56.79 42.075 -56.66 42.225)
MU9413/2/ix2031/2 U9413/2/ix2031/OUT U9413/2/ix2019/B U9413/2/ix2031/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-56.21 42.075 -56.08 42.225)
MU9413/2/ix2031/3 U9413/2/ix2031/3 wrData[28] U9413/2/ix2031/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-55.63 42.075 -55.5 42.225)
MU9413/2/ix2031/4 G_DG U9413/2/ix2019/D U9413/2/ix2031/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-55.05 42.075 -54.92 42.225)
MU9413/2/reg_r_shiftReg_29_/1 G_DG U9413/2/CLK U9413/2/35 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-71.115 42.075 -70.985 42.225)
MU9413/2/reg_r_shiftReg_29_/2 U9413/2/36 U9413/2/35 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-70.535 42.075 -70.405 42.225)
MU9413/2/reg_r_shiftReg_29_/3 U9413/2/reg_r_shiftReg_29_/4 U9413/2/ix397/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-69.445 42.075 -69.315 42.225)
MU9413/2/reg_r_shiftReg_29_/4 U9413/2/39 U9413/2/35 U9413/2/reg_r_shiftReg_29_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-68.93 42.075 -68.8 42.225)
MU9413/2/reg_r_shiftReg_29_/5 U9413/2/40 U9413/2/39 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-67.84 42.075 -67.71 42.225)
MU9413/2/reg_r_shiftReg_29_/6 U9413/2/reg_r_shiftReg_29_/7 U9413/2/CLB U9413/2/39 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-66.47 42.075 -66.34 42.225)
MU9413/2/reg_r_shiftReg_29_/7 U9413/2/reg_r_shiftReg_29_/8 U9413/2/40 U9413/2/reg_r_shiftReg_29_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-65.99 42.075 -65.86 42.225)
MU9413/2/reg_r_shiftReg_29_/8 G_DG U9413/2/36 U9413/2/reg_r_shiftReg_29_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-65.51 42.075 -65.38 42.225)
MU9413/2/reg_r_shiftReg_29_/9 U9413/2/reg_r_shiftReg_29_/9 U9413/2/40 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-64.42 42.075 -64.29 42.225)
MU9413/2/reg_r_shiftReg_29_/10 U9413/2/reg_r_shiftReg_29_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_29_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-63.91 42.075 -63.78 42.225)
MU9413/2/reg_r_shiftReg_29_/11 U9413/2/43 U9413/2/36 U9413/2/reg_r_shiftReg_29_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-63.49 42.075 -63.36 42.225)
MU9413/2/reg_r_shiftReg_29_/12 U9413/2/44 U9413/2/43 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-62.4 42.075 -62.27 42.225)
MU9413/2/reg_r_shiftReg_29_/13 U9413/2/45 U9413/2/35 U9413/2/43 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-61.04 42.075 -60.91 42.225)
MU9413/2/reg_r_shiftReg_29_/14 U9413/2/reg_r_shiftReg_29_/14 U9413/2/CLB U9413/2/45 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-60.46 42.075 -60.33 42.225)
MU9413/2/reg_r_shiftReg_29_/15 G_DG U9413/2/44 U9413/2/reg_r_shiftReg_29_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-60.15 42.075 -60.02 42.225)
MU9413/2/reg_r_shiftReg_29_/16 wrData[28] U9413/2/45 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-59.06 42.075 -58.93 42.225)
MU9413/2/reg_r_shiftReg_29_/17 U9413/2/reg_r_shiftReg_29_/QB U9413/2/44 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-57.97 42.075 -57.84 42.225)
MU9413/2/ix2025/1 U9413/2/ix2025/1 rdData[29] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-74.035 42.075 -73.905 42.225)
MU9413/2/ix2025/2 U9413/reg_r_shiftReg_47_\Cross U9413/2/ix2019/B U9413/2/ix2025/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-73.455 42.075 -73.325 42.225)
MU9413/2/ix2025/3 U9413/2/ix2025/3 wrData[29] U9413/reg_r_shiftReg_47_\Cross G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-72.875 42.075 -72.745 42.225)
MU9413/2/ix2025/4 G_DG U9413/2/ix2019/D U9413/2/ix2025/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-72.295 42.075 -72.165 42.225)
MU9413/2/ix2021/1 U9413/2/ix2021/1 wrData[29] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-75.795 42.075 -75.665 42.225)
MU9413/2/ix2021/2 U9413/2/ix2021/OUT U9413/2/ix2021/B U9413/2/ix2021/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-75.215 42.075 -75.085 42.225)
MU9413/2/ix2019/1 U9413/2/ix2019/1 rdData[30] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-78.715 42.075 -78.585 42.225)
MU9413/2/ix2019/2 U9413/2/ix2019/OUT U9413/2/ix2019/B U9413/2/ix2019/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-78.135 42.075 -78.005 42.225)
MU9413/2/ix2019/3 U9413/2/ix2019/3 wrData[30] U9413/2/ix2019/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-77.555 42.075 -77.425 42.225)
MU9413/2/ix2019/4 G_DG U9413/2/ix2019/D U9413/2/ix2019/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-76.975 42.075 -76.845 42.225)
MU9413/2/ix421/1 U9413/2/ix421/1 U9413/2/ix2019/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-80.475 42.075 -80.345 42.225)
MU9413/2/ix421/2 U9413/2/ix421/OUT U9413/2/ix2021/OUT U9413/2/ix421/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-79.895 42.075 -79.765 42.225)
MU9413/2/reg_r_shiftReg_31_/1 G_DG U9413/2/CLK U9413/2/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-94.8 42.075 -94.67 42.225)
MU9413/2/reg_r_shiftReg_31_/2 U9413/2/5 U9413/2/4 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-94.22 42.075 -94.09 42.225)
MU9413/2/reg_r_shiftReg_31_/3 U9413/2/reg_r_shiftReg_31_/4 U9413/2/ix421/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-93.13 42.075 -93 42.225)
MU9413/2/reg_r_shiftReg_31_/4 U9413/2/8 U9413/2/4 U9413/2/reg_r_shiftReg_31_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-92.615 42.075 -92.485 42.225)
MU9413/2/reg_r_shiftReg_31_/5 U9413/2/9 U9413/2/8 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-91.525 42.075 -91.395 42.225)
MU9413/2/reg_r_shiftReg_31_/6 U9413/2/reg_r_shiftReg_31_/7 U9413/2/CLB U9413/2/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-90.155 42.075 -90.025 42.225)
MU9413/2/reg_r_shiftReg_31_/7 U9413/2/reg_r_shiftReg_31_/8 U9413/2/9 U9413/2/reg_r_shiftReg_31_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-89.675 42.075 -89.545 42.225)
MU9413/2/reg_r_shiftReg_31_/8 G_DG U9413/2/5 U9413/2/reg_r_shiftReg_31_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-89.195 42.075 -89.065 42.225)
MU9413/2/reg_r_shiftReg_31_/9 U9413/2/reg_r_shiftReg_31_/9 U9413/2/9 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-88.105 42.075 -87.975 42.225)
MU9413/2/reg_r_shiftReg_31_/10 U9413/2/reg_r_shiftReg_31_/10 U9413/2/CLB U9413/2/reg_r_shiftReg_31_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-87.595 42.075 -87.465 42.225)
MU9413/2/reg_r_shiftReg_31_/11 U9413/2/12 U9413/2/5 U9413/2/reg_r_shiftReg_31_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-87.175 42.075 -87.045 42.225)
MU9413/2/reg_r_shiftReg_31_/12 U9413/2/13 U9413/2/12 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-86.085 42.075 -85.955 42.225)
MU9413/2/reg_r_shiftReg_31_/13 U9413/2/14 U9413/2/4 U9413/2/12 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-84.725 42.075 -84.595 42.225)
MU9413/2/reg_r_shiftReg_31_/14 U9413/2/reg_r_shiftReg_31_/14 U9413/2/CLB U9413/2/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-84.145 42.075 -84.015 42.225)
MU9413/2/reg_r_shiftReg_31_/15 G_DG U9413/2/13 U9413/2/reg_r_shiftReg_31_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-83.835 42.075 -83.705 42.225)
MU9413/2/reg_r_shiftReg_31_/16 wrData[30] U9413/2/14 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-82.745 42.075 -82.615 42.225)
MU9413/2/reg_r_shiftReg_31_/17 U9413/2/reg_r_shiftReg_31_/QB U9413/2/13 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-81.655 42.075 -81.525 42.225)
MU9413/3/1 G_DS CLK U9413/3/2 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-98.32 32.25 -98.19 32.55)
MU9413/3/2 U9413/3/CLK U9413/3/2 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-97.74 32.25 -97.61 32.55)
MU9413/3/3 G_DS CLK U9413/3/3 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-96.56 32.25 -96.43 32.55)
MU9413/3/4 U9413/3/CLK U9413/3/3 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-95.98 32.25 -95.85 32.55)
MU9413/3/5 G_DS U9413/SEL U9413/3/5 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-94.8 32.035 -94.67 32.335)
MU9413/3/6 U9413/3/6 U9413/3/5 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-94.22 32.035 -94.09 32.555)
MU9413/3/7 U9413/3/7 cmd[1] U9413/3/6 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-93.64 32.035 -93.51 32.555)
MU9413/3/8 U9413/3/9 cmd[2] U9413/3/7 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-93.06 32.035 -92.93 32.555)
MU9413/3/9 G_DS U9413/SEL U9413/3/9 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-92.48 32.035 -92.35 32.555)
MU9413/3/10 U9413/3/ix1846/OUT U9413/3/7 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-91.9 32.25 -91.77 32.55)
MU9413/3/11 G_DS U9413/3/CLK U9413/3/12 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-90.72 32.25 -90.59 32.55)
MU9413/3/12 U9413/3/13 U9413/3/12 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-90.14 32.25 -90.01 32.55)
MU9413/3/13 U9413/3/14 U9413/3/ix1846/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-89.05 32.25 -88.92 32.64)
MU9413/3/14 U9413/3/16 U9413/3/13 U9413/3/14 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-88.535 32.25 -88.405 32.64)
MU9413/3/15 U9413/3/17 U9413/3/16 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-87.445 32.25 -87.315 32.55)
MU9413/3/16 U9413/3/18 U9413/3/12 U9413/3/16 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-86.355 32.25 -86.225 32.64)
MU9413/3/17 G_DS U9413/3/CLB U9413/3/18 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-85.735 32.25 -85.605 32.64)
MU9413/3/18 U9413/3/18 U9413/3/17 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-85.115 32.25 -84.985 32.64)
MU9413/3/19 U9413/3/19 U9413/3/17 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-84.025 32.25 -83.895 32.64)
MU9413/3/20 U9413/3/20 U9413/3/12 U9413/3/19 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-83.715 32.25 -83.585 32.64)
MU9413/3/21 U9413/3/21 U9413/3/20 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-82.005 32.25 -81.875 32.55)
MU9413/3/22 U9413/3/22 U9413/3/13 U9413/3/20 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-80.915 32.25 -80.785 32.64)
MU9413/3/23 G_DS U9413/3/CLB U9413/3/22 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-80.335 32.25 -80.205 32.64)
MU9413/3/24 U9413/3/22 U9413/3/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-79.755 32.25 -79.625 32.55)
MU9413/3/25 cmd[2] U9413/3/22 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-78.665 32.25 -78.535 32.55)
MU9413/3/26 U9413/3/reg_r_shiftReg_47_/QB U9413/3/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-77.575 32.25 -77.445 32.55)
MU9413/3/27 U9413/3/25 rdData[31] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-76.395 32.035 -76.265 32.555)
MU9413/3/28 U9413/3/ix1993/OUT wrData[31] U9413/3/25 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-75.815 32.035 -75.685 32.555)
MU9413/3/29 U9413/3/25 U9413/2/ix2019/D U9413/3/ix1993/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-75.235 32.035 -75.105 32.555)
MU9413/3/30 G_DS U9413/2/ix2019/B U9413/3/25 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-74.655 32.035 -74.525 32.555)
MU9413/3/31 U9413/3/ix2015/OUT wrData[30] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-73.475 32.25 -73.345 32.51)
MU9413/3/32 G_DS U9413/2/ix2021/B U9413/3/ix2015/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-72.895 32.25 -72.765 32.51)
MU9413/3/33 U9413/3/ix433/OUT U9413/3/ix1993/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-71.715 32.25 -71.585 32.51)
MU9413/3/34 G_DS U9413/3/ix2015/OUT U9413/3/ix433/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-71.135 32.25 -71.005 32.51)
MU9413/3/35 U9413/3/ix2027/OUT wrData[28] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-69.955 32.25 -69.825 32.51)
MU9413/3/36 G_DS U9413/2/ix2021/B U9413/3/ix2027/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-69.375 32.25 -69.245 32.51)
MU9413/3/37 G_DS U9413/3/CLK U9413/3/40 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-68.195 32.25 -68.065 32.55)
MU9413/3/38 U9413/3/41 U9413/3/40 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-67.615 32.25 -67.485 32.55)
MU9413/3/39 U9413/3/42 U9413/3/ix433/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-66.525 32.25 -66.395 32.64)
MU9413/3/40 U9413/3/44 U9413/3/41 U9413/3/42 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-66.01 32.25 -65.88 32.64)
MU9413/3/41 U9413/3/45 U9413/3/44 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-64.92 32.25 -64.79 32.55)
MU9413/3/42 U9413/3/46 U9413/3/40 U9413/3/44 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-63.83 32.25 -63.7 32.64)
MU9413/3/43 G_DS U9413/3/CLB U9413/3/46 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-63.21 32.25 -63.08 32.64)
MU9413/3/44 U9413/3/46 U9413/3/45 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-62.59 32.25 -62.46 32.64)
MU9413/3/45 U9413/3/47 U9413/3/45 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-61.5 32.25 -61.37 32.64)
MU9413/3/46 U9413/3/48 U9413/3/40 U9413/3/47 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-61.19 32.25 -61.06 32.64)
MU9413/3/47 U9413/3/49 U9413/3/48 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-59.48 32.25 -59.35 32.55)
MU9413/3/48 U9413/3/50 U9413/3/41 U9413/3/48 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-58.39 32.25 -58.26 32.64)
MU9413/3/49 G_DS U9413/3/CLB U9413/3/50 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-57.81 32.25 -57.68 32.64)
MU9413/3/50 U9413/3/50 U9413/3/49 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-57.23 32.25 -57.1 32.55)
MU9413/3/51 wrData[31] U9413/3/50 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-56.14 32.25 -56.01 32.55)
MU9413/3/52 U9413/3/reg_r_shiftReg_32_/QB U9413/3/49 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-55.05 32.25 -54.92 32.55)
MU9413/3/53 U9413/3/53 rdData[27] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-53.87 32.035 -53.74 32.555)
MU9413/3/54 U9413/3/ix2037/OUT wrData[27] U9413/3/53 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-53.29 32.035 -53.16 32.555)
MU9413/3/55 U9413/3/53 U9413/2/ix2019/D U9413/3/ix2037/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-52.71 32.035 -52.58 32.555)
MU9413/3/56 G_DS U9413/2/ix2019/B U9413/3/53 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-52.13 32.035 -52 32.555)
MU9413/3/57 U9413/3/ix385/OUT U9413/3/ix2037/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-50.95 32.25 -50.82 32.51)
MU9413/3/58 G_DS U9413/3/ix2039/OUT U9413/3/ix385/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-50.37 32.25 -50.24 32.51)
MU9413/3/59 U9413/3/ix2039/OUT wrData[26] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-49.19 32.25 -49.06 32.51)
MU9413/3/60 G_DS U9413/2/ix2045/B U9413/3/ix2039/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-48.61 32.25 -48.48 32.51)
MU9413/3/61 G_DS U9413/3/CLK U9413/3/65 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-47.43 32.25 -47.3 32.55)
MU9413/3/62 U9413/3/66 U9413/3/65 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-46.85 32.25 -46.72 32.55)
MU9413/3/63 U9413/3/67 U9413/2/ix373/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-45.76 32.25 -45.63 32.64)
MU9413/3/64 U9413/3/69 U9413/3/66 U9413/3/67 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-45.245 32.25 -45.115 32.64)
MU9413/3/65 U9413/3/70 U9413/3/69 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-44.155 32.25 -44.025 32.55)
MU9413/3/66 U9413/3/71 U9413/3/65 U9413/3/69 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-43.065 32.25 -42.935 32.64)
MU9413/3/67 G_DS U9413/3/CLB U9413/3/71 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-42.445 32.25 -42.315 32.64)
MU9413/3/68 U9413/3/71 U9413/3/70 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-41.825 32.25 -41.695 32.64)
MU9413/3/69 U9413/3/72 U9413/3/70 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-40.735 32.25 -40.605 32.64)
MU9413/3/70 U9413/3/73 U9413/3/65 U9413/3/72 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-40.425 32.25 -40.295 32.64)
MU9413/3/71 U9413/3/74 U9413/3/73 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-38.715 32.25 -38.585 32.55)
MU9413/3/72 U9413/3/75 U9413/3/66 U9413/3/73 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-37.625 32.25 -37.495 32.64)
MU9413/3/73 G_DS U9413/3/CLB U9413/3/75 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-37.045 32.25 -36.915 32.64)
MU9413/3/74 U9413/3/75 U9413/3/74 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-36.465 32.25 -36.335 32.55)
MU9413/3/75 wrData[26] U9413/3/75 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-35.375 32.25 -35.245 32.55)
MU9413/3/76 U9413/3/reg_r_shiftReg_27_/QB U9413/3/74 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-34.285 32.25 -34.155 32.55)
MU9413/3/77 U9413/3/78 rdData[24] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-33.105 32.035 -32.975 32.555)
MU9413/3/78 U9413/3/ix2055/OUT wrData[24] U9413/3/78 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-32.525 32.035 -32.395 32.555)
MU9413/3/79 U9413/3/78 U9413/2/ix2019/D U9413/3/ix2055/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-31.945 32.035 -31.815 32.555)
MU9413/3/80 G_DS U9413/2/ix2019/B U9413/3/78 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-31.365 32.035 -31.235 32.555)
MU9413/3/81 U9413/3/ix349/OUT U9413/3/ix2055/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-30.185 32.25 -30.055 32.51)
MU9413/3/82 G_DS U9413/3/ix2057/OUT U9413/3/ix349/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-29.605 32.25 -29.475 32.51)
MU9413/3/83 U9413/3/ix2057/OUT wrData[23] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-28.425 32.25 -28.295 32.51)
MU9413/3/84 G_DS U9413/2/ix2045/B U9413/3/ix2057/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-27.845 32.25 -27.715 32.51)
MU9413/3/85 U9413/3/ix2063/OUT wrData[22] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-26.665 32.25 -26.535 32.51)
MU9413/3/86 G_DS U9413/2/ix2045/B U9413/3/ix2063/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-26.085 32.25 -25.955 32.51)
MU9413/3/87 U9413/3/ix337/OUT U9413/2/ix2061/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-24.905 32.25 -24.775 32.51)
MU9413/3/88 G_DS U9413/3/ix2063/OUT U9413/3/ix337/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-24.325 32.25 -24.195 32.51)
MU9413/3/89 G_DS U9413/3/CLK U9413/3/96 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-23.145 32.25 -23.015 32.55)
MU9413/3/90 U9413/3/97 U9413/3/96 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-22.565 32.25 -22.435 32.55)
MU9413/3/91 U9413/3/98 U9413/3/ix337/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-21.475 32.25 -21.345 32.64)
MU9413/3/92 U9413/3/100 U9413/3/97 U9413/3/98 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-20.96 32.25 -20.83 32.64)
MU9413/3/93 U9413/3/101 U9413/3/100 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-19.87 32.25 -19.74 32.55)
MU9413/3/94 U9413/3/102 U9413/3/96 U9413/3/100 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-18.78 32.25 -18.65 32.64)
MU9413/3/95 G_DS U9413/3/CLB U9413/3/102 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-18.16 32.25 -18.03 32.64)
MU9413/3/96 U9413/3/102 U9413/3/101 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-17.54 32.25 -17.41 32.64)
MU9413/3/97 U9413/3/103 U9413/3/101 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-16.45 32.25 -16.32 32.64)
MU9413/3/98 U9413/3/104 U9413/3/96 U9413/3/103 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-16.14 32.25 -16.01 32.64)
MU9413/3/99 U9413/3/105 U9413/3/104 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-14.43 32.25 -14.3 32.55)
MU9413/3/100 U9413/3/106 U9413/3/97 U9413/3/104 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-13.34 32.25 -13.21 32.64)
MU9413/3/101 G_DS U9413/3/CLB U9413/3/106 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-12.76 32.25 -12.63 32.64)
MU9413/3/102 U9413/3/106 U9413/3/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-12.18 32.25 -12.05 32.55)
MU9413/3/103 wrData[23] U9413/3/106 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-11.09 32.25 -10.96 32.55)
MU9413/3/104 U9413/3/reg_r_shiftReg_24_/QB U9413/3/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-10 32.25 -9.87 32.55)
MU9413/3/105 U9413/3/109 rdData[21] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(-8.82 32.035 -8.69 32.555)
MU9413/3/106 U9413/3/ix2073/OUT wrData[21] U9413/3/109 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-8.24 32.035 -8.11 32.555)
MU9413/3/107 U9413/3/109 U9413/2/ix2067/D U9413/3/ix2073/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(-7.66 32.035 -7.53 32.555)
MU9413/3/108 G_DS U9413/2/ix2067/B U9413/3/109 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(-7.08 32.035 -6.95 32.555)
MU9413/3/109 G_DS U9413/3/CLK U9413/3/115 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-5.9 32.25 -5.77 32.55)
MU9413/3/110 U9413/3/116 U9413/3/115 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-5.32 32.25 -5.19 32.55)
MU9413/3/111 U9413/3/117 U9413/3/ix301/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-4.23 32.25 -4.1 32.64)
MU9413/3/112 U9413/3/119 U9413/3/116 U9413/3/117 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-3.715 32.25 -3.585 32.64)
MU9413/3/113 U9413/3/120 U9413/3/119 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-2.625 32.25 -2.495 32.55)
MU9413/3/114 U9413/3/121 U9413/3/115 U9413/3/119 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-1.535 32.25 -1.405 32.64)
MU9413/3/115 G_DS U9413/3/CLB U9413/3/121 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-0.915 32.25 -0.785 32.64)
MU9413/3/116 U9413/3/121 U9413/3/120 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-0.295 32.25 -0.165 32.64)
MU9413/3/117 U9413/3/122 U9413/3/120 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(0.795 32.25 0.925 32.64)
MU9413/3/118 U9413/3/123 U9413/3/115 U9413/3/122 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(1.105 32.25 1.235 32.64)
MU9413/3/119 U9413/3/124 U9413/3/123 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(2.815 32.25 2.945 32.55)
MU9413/3/120 U9413/3/125 U9413/3/116 U9413/3/123 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(3.905 32.25 4.035 32.64)
MU9413/3/121 G_DS U9413/3/CLB U9413/3/125 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(4.485 32.25 4.615 32.64)
MU9413/3/122 U9413/3/125 U9413/3/124 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(5.065 32.25 5.195 32.55)
MU9413/3/123 wrData[20] U9413/3/125 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(6.155 32.25 6.285 32.55)
MU9413/3/124 U9413/3/reg_r_shiftReg_21_/QB U9413/3/124 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(7.245 32.25 7.375 32.55)
MU9413/3/125 U9413/3/ix301/OUT U9413/2/ix2079/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(8.425 32.25 8.555 32.51)
MU9413/3/126 G_DS U9413/3/ix2081/OUT U9413/3/ix301/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(9.005 32.25 9.135 32.51)
MU9413/3/127 U9413/3/ix2081/OUT wrData[19] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(10.185 32.25 10.315 32.51)
MU9413/3/128 G_DS U9413/2/ix2045/B U9413/3/ix2081/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(10.765 32.25 10.895 32.51)
MU9413/3/129 G_DS U9413/3/ix2292/A U9413/3/135 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(11.945 32.25 12.075 32.55)
MU9413/3/130 U9413/2/ix2067/B U9413/3/135 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(12.525 32.25 12.655 32.55)
MU9413/3/131 U9413/3/137 rdData[17] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(13.705 32.035 13.835 32.555)
MU9413/3/132 U9413/3/ix2097/OUT wrData[17] U9413/3/137 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(14.285 32.035 14.415 32.555)
MU9413/3/133 U9413/3/137 U9413/2/ix2067/D U9413/3/ix2097/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(14.865 32.035 14.995 32.555)
MU9413/3/134 G_DS U9413/2/ix2067/B U9413/3/137 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(15.445 32.035 15.575 32.555)
MU9413/3/135 G_DS U9413/3/CLK U9413/3/143 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(16.625 32.25 16.755 32.55)
MU9413/3/136 U9413/3/144 U9413/3/143 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(17.205 32.25 17.335 32.55)
MU9413/3/137 U9413/3/145 U9413/2/ix289/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(18.295 32.25 18.425 32.64)
MU9413/3/138 U9413/3/147 U9413/3/144 U9413/3/145 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(18.81 32.25 18.94 32.64)
MU9413/3/139 U9413/3/148 U9413/3/147 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(19.9 32.25 20.03 32.55)
MU9413/3/140 U9413/3/149 U9413/3/143 U9413/3/147 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(20.99 32.25 21.12 32.64)
MU9413/3/141 G_DS U9413/3/CLB U9413/3/149 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(21.61 32.25 21.74 32.64)
MU9413/3/142 U9413/3/149 U9413/3/148 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(22.23 32.25 22.36 32.64)
MU9413/3/143 U9413/3/150 U9413/3/148 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(23.32 32.25 23.45 32.64)
MU9413/3/144 U9413/3/151 U9413/3/143 U9413/3/150 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(23.63 32.25 23.76 32.64)
MU9413/3/145 U9413/3/152 U9413/3/151 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(25.34 32.25 25.47 32.55)
MU9413/3/146 U9413/3/153 U9413/3/144 U9413/3/151 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(26.43 32.25 26.56 32.64)
MU9413/3/147 G_DS U9413/3/CLB U9413/3/153 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(27.01 32.25 27.14 32.64)
MU9413/3/148 U9413/3/153 U9413/3/152 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(27.59 32.25 27.72 32.55)
MU9413/3/149 wrData[19] U9413/3/153 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(28.68 32.25 28.81 32.55)
MU9413/3/150 U9413/3/reg_r_shiftReg_20_/QB U9413/3/152 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(29.77 32.25 29.9 32.55)
MU9413/3/151 U9413/3/156 rdData[16] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(30.95 32.035 31.08 32.555)
MU9413/3/152 U9413/3/ix2103/OUT wrData[16] U9413/3/156 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(31.53 32.035 31.66 32.555)
MU9413/3/153 U9413/3/156 U9413/2/ix2067/D U9413/3/ix2103/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(32.11 32.035 32.24 32.555)
MU9413/3/154 G_DS U9413/2/ix2067/B U9413/3/156 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(32.69 32.035 32.82 32.555)
MU9413/3/155 U9413/3/162 rdData[14] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(33.87 32.035 34 32.555)
MU9413/3/156 U9413/3/ix2115/OUT wrData[14] U9413/3/162 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(34.45 32.035 34.58 32.555)
MU9413/3/157 U9413/3/162 U9413/2/ix2067/D U9413/3/ix2115/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(35.03 32.035 35.16 32.555)
MU9413/3/158 G_DS U9413/2/ix2067/B U9413/3/162 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(35.61 32.035 35.74 32.555)
MU9413/3/159 U9413/3/ix253/OUT U9413/3/ix2103/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(36.79 32.25 36.92 32.51)
MU9413/3/160 G_DS U9413/2/ix2105/OUT U9413/3/ix253/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(37.37 32.25 37.5 32.51)
MU9413/3/161 G_DS U9413/3/CLK U9413/3/171 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(38.55 32.25 38.68 32.55)
MU9413/3/162 U9413/3/172 U9413/3/171 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(39.13 32.25 39.26 32.55)
MU9413/3/163 U9413/3/173 U9413/3/ix253/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(40.22 32.25 40.35 32.64)
MU9413/3/164 U9413/3/175 U9413/3/172 U9413/3/173 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(40.735 32.25 40.865 32.64)
MU9413/3/165 U9413/3/176 U9413/3/175 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(41.825 32.25 41.955 32.55)
MU9413/3/166 U9413/3/177 U9413/3/171 U9413/3/175 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(42.915 32.25 43.045 32.64)
MU9413/3/167 G_DS U9413/3/CLB U9413/3/177 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(43.535 32.25 43.665 32.64)
MU9413/3/168 U9413/3/177 U9413/3/176 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(44.155 32.25 44.285 32.64)
MU9413/3/169 U9413/3/178 U9413/3/176 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(45.245 32.25 45.375 32.64)
MU9413/3/170 U9413/3/179 U9413/3/171 U9413/3/178 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(45.555 32.25 45.685 32.64)
MU9413/3/171 U9413/3/180 U9413/3/179 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(47.265 32.25 47.395 32.55)
MU9413/3/172 U9413/3/181 U9413/3/172 U9413/3/179 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(48.355 32.25 48.485 32.64)
MU9413/3/173 G_DS U9413/3/CLB U9413/3/181 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(48.935 32.25 49.065 32.64)
MU9413/3/174 U9413/3/181 U9413/3/180 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(49.515 32.25 49.645 32.55)
MU9413/3/175 wrData[16] U9413/3/181 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(50.605 32.25 50.735 32.55)
MU9413/3/176 U9413/3/reg_r_shiftReg_17_/QB U9413/3/180 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(51.695 32.25 51.825 32.55)
MU9413/3/177 U9413/3/ix217/OUT U9413/2/ix2121/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(52.875 32.25 53.005 32.51)
MU9413/3/178 G_DS U9413/3/ix2123/OUT U9413/3/ix217/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(53.455 32.25 53.585 32.51)
MU9413/3/179 U9413/3/ix2123/OUT wrData[12] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(54.635 32.25 54.765 32.51)
MU9413/3/180 G_DS U9413/2/ix2093/B U9413/3/ix2123/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(55.215 32.25 55.345 32.51)
MU9413/3/181 G_DS U9413/3/ix2292/A U9413/3/191 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(56.395 32.25 56.525 32.55)
MU9413/3/182 U9413/2/ix2121/B U9413/3/191 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(56.975 32.25 57.105 32.55)
MU9413/3/183 U9413/3/ix193/OUT U9413/2/ix2133/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(58.155 32.25 58.285 32.51)
MU9413/3/184 G_DS U9413/3/ix193/B U9413/3/ix193/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(58.735 32.25 58.865 32.51)
MU9413/3/185 U9413/3/ix193/B wrData[10] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(59.915 32.25 60.045 32.51)
MU9413/3/186 G_DS U9413/2/ix2093/B U9413/3/ix193/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(60.495 32.25 60.625 32.51)
MU9413/3/187 G_DS U9413/3/CLK U9413/3/199 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(61.675 32.25 61.805 32.55)
MU9413/3/188 U9413/3/200 U9413/3/199 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(62.255 32.25 62.385 32.55)
MU9413/3/189 U9413/3/201 U9413/2/ix181/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(63.345 32.25 63.475 32.64)
MU9413/3/190 U9413/3/203 U9413/3/200 U9413/3/201 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(63.86 32.25 63.99 32.64)
MU9413/3/191 U9413/3/204 U9413/3/203 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(64.95 32.25 65.08 32.55)
MU9413/3/192 U9413/3/205 U9413/3/199 U9413/3/203 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(66.04 32.25 66.17 32.64)
MU9413/3/193 G_DS U9413/3/CLB U9413/3/205 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(66.66 32.25 66.79 32.64)
MU9413/3/194 U9413/3/205 U9413/3/204 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(67.28 32.25 67.41 32.64)
MU9413/3/195 U9413/3/206 U9413/3/204 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(68.37 32.25 68.5 32.64)
MU9413/3/196 U9413/3/207 U9413/3/199 U9413/3/206 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(68.68 32.25 68.81 32.64)
MU9413/3/197 U9413/3/208 U9413/3/207 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(70.39 32.25 70.52 32.55)
MU9413/3/198 U9413/3/209 U9413/3/200 U9413/3/207 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(71.48 32.25 71.61 32.64)
MU9413/3/199 G_DS U9413/3/CLB U9413/3/209 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(72.06 32.25 72.19 32.64)
MU9413/3/200 U9413/3/209 U9413/3/208 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(72.64 32.25 72.77 32.55)
MU9413/3/201 wrData[10] U9413/3/209 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(73.73 32.25 73.86 32.55)
MU9413/3/202 U9413/3/reg_r_shiftReg_11_/QB U9413/3/208 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(74.82 32.25 74.95 32.55)
MU9413/3/203 U9413/3/212 rdData[8] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(76 32.035 76.13 32.555)
MU9413/3/204 U9413/3/ix2151/OUT wrData[8] U9413/3/212 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(76.58 32.035 76.71 32.555)
MU9413/3/205 U9413/3/212 U9413/2/ix2121/D U9413/3/ix2151/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(77.16 32.035 77.29 32.555)
MU9413/3/206 G_DS U9413/2/ix2121/B U9413/3/212 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(77.74 32.035 77.87 32.555)
MU9413/3/207 U9413/3/218 rdData[7] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(78.92 32.035 79.05 32.555)
MU9413/3/208 U9413/3/ix2157/OUT wrData[7] U9413/3/218 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(79.5 32.035 79.63 32.555)
MU9413/3/209 U9413/3/218 U9413/2/ix2121/D U9413/3/ix2157/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(80.08 32.035 80.21 32.555)
MU9413/3/210 G_DS U9413/2/ix2121/B U9413/3/218 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(80.66 32.035 80.79 32.555)
MU9413/3/211 G_DS U9413/3/ix2292/A U9413/3/225 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(81.84 32.25 81.97 32.55)
MU9413/3/212 U9413/2/ix1948/B U9413/3/225 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(82.42 32.25 82.55 32.55)
MU9413/3/213 U9413/3/ix133/OUT U9413/3/ix133/A G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(83.6 32.25 83.73 32.51)
MU9413/3/214 G_DS U9413/3/ix133/B U9413/3/ix133/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(84.18 32.25 84.31 32.51)
MU9413/3/215 U9413/3/230 rdData[6] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(85.36 32.035 85.49 32.555)
MU9413/3/216 U9413/3/ix133/A wrData[6] U9413/3/230 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(85.94 32.035 86.07 32.555)
MU9413/3/217 U9413/3/230 U9413/2/ix2121/D U9413/3/ix133/A G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(86.52 32.035 86.65 32.555)
MU9413/3/218 G_DS U9413/2/ix2121/B U9413/3/230 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(87.1 32.035 87.23 32.555)
MU9413/3/219 U9413/3/ix133/B wrData[5] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(88.28 32.25 88.41 32.51)
MU9413/3/220 G_DS U9413/2/ix2147/B U9413/3/ix133/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(88.86 32.25 88.99 32.51)
MU9413/3/221 G_DS U9413/3/CLK U9413/3/239 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(90.04 32.25 90.17 32.55)
MU9413/3/222 U9413/3/240 U9413/3/239 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(90.62 32.25 90.75 32.55)
MU9413/3/223 U9413/3/241 U9413/3/ix109/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(91.71 32.25 91.84 32.64)
MU9413/3/224 U9413/3/243 U9413/3/240 U9413/3/241 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(92.225 32.25 92.355 32.64)
MU9413/3/225 U9413/3/244 U9413/3/243 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(93.315 32.25 93.445 32.55)
MU9413/3/226 U9413/3/245 U9413/3/239 U9413/3/243 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(94.405 32.25 94.535 32.64)
MU9413/3/227 G_DS U9413/3/CLB U9413/3/245 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(95.025 32.25 95.155 32.64)
MU9413/3/228 U9413/3/245 U9413/3/244 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(95.645 32.25 95.775 32.64)
MU9413/3/229 U9413/3/246 U9413/3/244 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(96.735 32.25 96.865 32.64)
MU9413/3/230 U9413/3/247 U9413/3/239 U9413/3/246 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(97.045 32.25 97.175 32.64)
MU9413/3/231 U9413/3/248 U9413/3/247 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(98.755 32.25 98.885 32.55)
MU9413/3/232 U9413/3/249 U9413/3/240 U9413/3/247 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(99.845 32.25 99.975 32.64)
MU9413/3/233 G_DS U9413/3/CLB U9413/3/249 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(100.425 32.25 100.555 32.64)
MU9413/3/234 U9413/3/249 U9413/3/248 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(101.005 32.25 101.135 32.55)
MU9413/3/235 wrData[4] U9413/3/249 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(102.095 32.25 102.225 32.55)
MU9413/3/236 U9413/3/reg_r_shiftReg_5_/QB U9413/3/248 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(103.185 32.25 103.315 32.55)
MU9413/3/237 U9413/3/ix109/OUT U9413/2/ix2175/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(104.365 32.25 104.495 32.51)
MU9413/3/238 G_DS U9413/3/ix109/B U9413/3/ix109/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(104.945 32.25 105.075 32.51)
MU9413/3/239 U9413/3/ix109/B wrData[3] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(106.125 32.25 106.255 32.51)
MU9413/3/240 G_DS U9413/2/ix2147/B U9413/3/ix109/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(106.705 32.25 106.835 32.51)
MU9413/3/241 U9413/3/258 rdData[3] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(107.885 32.035 108.015 32.555)
MU9413/3/242 U9413/3/ix2181/OUT wrData[3] U9413/3/258 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(108.465 32.035 108.595 32.555)
MU9413/3/243 U9413/3/258 U9413/D U9413/3/ix2181/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(109.045 32.035 109.175 32.555)
MU9413/3/244 G_DS U9413/2/ix1948/B U9413/3/258 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(109.625 32.035 109.755 32.555)
MU9413/3/245 U9413/ix1786\Cross U9413/3/ix2187/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(110.805 32.25 110.935 32.51)
MU9413/3/246 G_DS U9413/2/ix2189/OUT U9413/ix1786\Cross G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(111.385 32.25 111.515 32.51)
MU9413/3/247 U9413/3/267 rdData[2] G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.35e-013 pd=1.09e-006 ps=2.03e-006 nrd=0.49926 nrs=0.85429  $(112.565 32.035 112.695 32.555)
MU9413/3/248 U9413/3/ix2187/OUT wrData[2] U9413/3/267 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(113.145 32.035 113.275 32.555)
MU9413/3/249 U9413/3/267 U9413/D U9413/3/ix2187/OUT G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.35e-013 pd=1.09e-006 ps=1.09e-006 nrd=0.49926 nrs=0.49926  $(113.725 32.035 113.855 32.555)
MU9413/3/250 G_DS U9413/2/ix1948/B U9413/3/267 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=2.31e-013 pd=2.03e-006 ps=1.09e-006 nrd=0.85429 nrs=0.49926  $(114.305 32.035 114.435 32.555)
MU9413/3/251 G_DS U9413/3/CLK U9413/3/271 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(115.485 32.25 115.615 32.55)
MU9413/3/252 U9413/3/272 U9413/3/271 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(116.065 32.25 116.195 32.55)
MU9413/3/253 U9413/3/273 U9413/3/ix1816/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(117.155 32.25 117.285 32.64)
MU9413/3/254 U9413/3/275 U9413/3/272 U9413/3/273 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(117.67 32.25 117.8 32.64)
MU9413/3/255 U9413/3/276 U9413/3/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(118.76 32.25 118.89 32.55)
MU9413/3/256 U9413/3/277 U9413/3/271 U9413/3/275 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(119.85 32.25 119.98 32.64)
MU9413/3/257 G_DS U9413/3/CLB U9413/3/277 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(120.47 32.25 120.6 32.64)
MU9413/3/258 U9413/3/277 U9413/3/276 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(121.09 32.25 121.22 32.64)
MU9413/3/259 U9413/3/278 U9413/3/276 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(122.18 32.25 122.31 32.64)
MU9413/3/260 U9413/3/279 U9413/3/271 U9413/3/278 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(122.49 32.25 122.62 32.64)
MU9413/3/261 U9413/3/280 U9413/3/279 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(124.2 32.25 124.33 32.55)
MU9413/3/262 U9413/3/281 U9413/3/272 U9413/3/279 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(125.29 32.25 125.42 32.64)
MU9413/3/263 G_DS U9413/3/CLB U9413/3/281 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(125.87 32.25 126 32.64)
MU9413/3/264 U9413/3/281 U9413/3/280 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(126.45 32.25 126.58 32.55)
MU9413/3/265 addr[11] U9413/3/281 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(127.54 32.25 127.67 32.55)
MU9413/3/266 U9413/3/reg_r_shiftReg_44_/QB U9413/3/280 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(128.63 32.25 128.76 32.55)
MU9413/3/267 G_DS U9413/SEL U9413/3/285 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(129.81 32.035 129.94 32.335)
MU9413/3/268 U9413/3/286 U9413/3/285 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(130.39 32.035 130.52 32.555)
MU9413/3/269 U9413/3/287 addr[10] U9413/3/286 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(130.97 32.035 131.1 32.555)
MU9413/3/270 U9413/3/289 addr[11] U9413/3/287 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(131.55 32.035 131.68 32.555)
MU9413/3/271 G_DS U9413/SEL U9413/3/289 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(132.13 32.035 132.26 32.555)
MU9413/3/272 U9413/3/ix1816/OUT U9413/3/287 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(132.71 32.25 132.84 32.55)
MU9413/3/273 G_DS U9413/SEL U9413/3/292 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(133.89 32.035 134.02 32.335)
MU9413/3/274 U9413/3/293 U9413/3/292 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(134.47 32.035 134.6 32.555)
MU9413/3/275 U9413/3/294 addr[9] U9413/3/293 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(135.05 32.035 135.18 32.555)
MU9413/3/276 U9413/3/295 addr[10] U9413/3/294 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(135.63 32.035 135.76 32.555)
MU9413/3/277 G_DS U9413/SEL U9413/3/295 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(136.21 32.035 136.34 32.555)
MU9413/3/278 U9413/3/DATA U9413/3/294 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(136.79 32.25 136.92 32.55)
MU9413/3/279 G_DS U9413/3/CLK U9413/3/296 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(137.97 32.25 138.1 32.55)
MU9413/3/280 U9413/3/297 U9413/3/296 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(138.55 32.25 138.68 32.55)
MU9413/3/281 U9413/3/298 U9413/3/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(139.64 32.25 139.77 32.64)
MU9413/3/282 U9413/3/299 U9413/3/297 U9413/3/298 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(140.155 32.25 140.285 32.64)
MU9413/3/283 U9413/3/300 U9413/3/299 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(141.245 32.25 141.375 32.55)
MU9413/3/284 U9413/3/301 U9413/3/296 U9413/3/299 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(142.335 32.25 142.465 32.64)
MU9413/3/285 G_DS U9413/3/CLB U9413/3/301 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(142.955 32.25 143.085 32.64)
MU9413/3/286 U9413/3/301 U9413/3/300 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(143.575 32.25 143.705 32.64)
MU9413/3/287 U9413/3/302 U9413/3/300 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(144.665 32.25 144.795 32.64)
MU9413/3/288 U9413/3/303 U9413/3/296 U9413/3/302 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(144.975 32.25 145.105 32.64)
MU9413/3/289 U9413/3/304 U9413/3/303 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(146.685 32.25 146.815 32.55)
MU9413/3/290 U9413/3/305 U9413/3/297 U9413/3/303 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(147.775 32.25 147.905 32.64)
MU9413/3/291 G_DS U9413/3/CLB U9413/3/305 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(148.355 32.25 148.485 32.64)
MU9413/3/292 U9413/3/305 U9413/3/304 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(148.935 32.25 149.065 32.55)
MU9413/3/293 addr[10] U9413/3/305 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(150.025 32.25 150.155 32.55)
MU9413/3/294 U9413/3/reg_r_shiftReg_43_/QB U9413/3/304 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(151.115 32.25 151.245 32.55)
MU9413/3/295 G_DS RST U9413/3/307 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(152.295 32.25 152.425 32.55)
MU9413/3/296 U9413/3/CLB U9413/3/307 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(152.875 32.25 153.005 32.55)
MU9413/3/297 G_DS RST U9413/3/308 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(154.055 32.25 154.185 32.55)
MU9413/3/298 U9413/3/CLB U9413/3/308 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(154.635 32.25 154.765 32.55)
MU9413/3/right_41/1 G_DG RST U9413/3/307 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(152.295 30.52 152.425 30.67)
MU9413/3/right_41/2 U9413/3/CLB U9413/3/307 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(152.875 30.52 153.005 30.67)
MU9413/3/right_40/1 G_DG RST U9413/3/308 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(154.055 30.52 154.185 30.67)
MU9413/3/right_40/2 U9413/3/CLB U9413/3/308 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(154.635 30.52 154.765 30.67)
MU9413/3/left_41/1 G_DG CLK U9413/3/2 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-98.32 30.52 -98.19 30.67)
MU9413/3/left_41/2 U9413/3/CLK U9413/3/2 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-97.74 30.52 -97.61 30.67)
MU9413/3/left_40/1 G_DG CLK U9413/3/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-96.56 30.52 -96.43 30.67)
MU9413/3/left_40/2 U9413/3/CLK U9413/3/3 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-95.98 30.52 -95.85 30.67)
MU9413/3/reg_r_shiftReg_43_/1 G_DG U9413/3/CLK U9413/3/296 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(137.97 30.52 138.1 30.67)
MU9413/3/reg_r_shiftReg_43_/2 U9413/3/297 U9413/3/296 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(138.55 30.52 138.68 30.67)
MU9413/3/reg_r_shiftReg_43_/3 U9413/3/reg_r_shiftReg_43_/4 U9413/3/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(139.64 30.52 139.77 30.67)
MU9413/3/reg_r_shiftReg_43_/4 U9413/3/299 U9413/3/296 U9413/3/reg_r_shiftReg_43_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(140.155 30.52 140.285 30.67)
MU9413/3/reg_r_shiftReg_43_/5 U9413/3/300 U9413/3/299 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(141.245 30.52 141.375 30.67)
MU9413/3/reg_r_shiftReg_43_/6 U9413/3/reg_r_shiftReg_43_/7 U9413/3/CLB U9413/3/299 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(142.615 30.52 142.745 30.67)
MU9413/3/reg_r_shiftReg_43_/7 U9413/3/reg_r_shiftReg_43_/8 U9413/3/300 U9413/3/reg_r_shiftReg_43_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(143.095 30.52 143.225 30.67)
MU9413/3/reg_r_shiftReg_43_/8 G_DG U9413/3/297 U9413/3/reg_r_shiftReg_43_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(143.575 30.52 143.705 30.67)
MU9413/3/reg_r_shiftReg_43_/9 U9413/3/reg_r_shiftReg_43_/9 U9413/3/300 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(144.665 30.52 144.795 30.67)
MU9413/3/reg_r_shiftReg_43_/10 U9413/3/reg_r_shiftReg_43_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_43_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(145.175 30.52 145.305 30.67)
MU9413/3/reg_r_shiftReg_43_/11 U9413/3/303 U9413/3/297 U9413/3/reg_r_shiftReg_43_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(145.595 30.52 145.725 30.67)
MU9413/3/reg_r_shiftReg_43_/12 U9413/3/304 U9413/3/303 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(146.685 30.52 146.815 30.67)
MU9413/3/reg_r_shiftReg_43_/13 U9413/3/305 U9413/3/296 U9413/3/303 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(148.045 30.52 148.175 30.67)
MU9413/3/reg_r_shiftReg_43_/14 U9413/3/reg_r_shiftReg_43_/14 U9413/3/CLB U9413/3/305 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(148.625 30.52 148.755 30.67)
MU9413/3/reg_r_shiftReg_43_/15 G_DG U9413/3/304 U9413/3/reg_r_shiftReg_43_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(148.935 30.52 149.065 30.67)
MU9413/3/reg_r_shiftReg_43_/16 addr[10] U9413/3/305 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(150.025 30.52 150.155 30.67)
MU9413/3/reg_r_shiftReg_43_/17 U9413/3/reg_r_shiftReg_43_/QB U9413/3/304 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(151.115 30.52 151.245 30.67)
MU9413/3/ix1806/1 G_DG U9413/SEL U9413/3/292 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(133.89 30.52 134.02 30.67)
MU9413/3/ix1806/2 U9413/3/ix1806/3 U9413/3/292 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(134.47 30.52 134.6 30.67)
MU9413/3/ix1806/3 U9413/3/294 addr[10] U9413/3/ix1806/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(135.05 30.52 135.18 30.67)
MU9413/3/ix1806/4 U9413/3/ix1806/5 addr[9] U9413/3/294 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(135.63 30.52 135.76 30.67)
MU9413/3/ix1806/5 G_DG U9413/SEL U9413/3/ix1806/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(136.21 30.52 136.34 30.67)
MU9413/3/ix1806/6 U9413/3/DATA U9413/3/294 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(136.79 30.52 136.92 30.67)
MU9413/3/ix1816/1 G_DG U9413/SEL U9413/3/285 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(129.81 30.52 129.94 30.67)
MU9413/3/ix1816/2 U9413/3/ix1816/3 U9413/3/285 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(130.39 30.52 130.52 30.67)
MU9413/3/ix1816/3 U9413/3/287 addr[11] U9413/3/ix1816/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(130.97 30.52 131.1 30.67)
MU9413/3/ix1816/4 U9413/3/ix1816/5 addr[10] U9413/3/287 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(131.55 30.52 131.68 30.67)
MU9413/3/ix1816/5 G_DG U9413/SEL U9413/3/ix1816/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(132.13 30.52 132.26 30.67)
MU9413/3/ix1816/6 U9413/3/ix1816/OUT U9413/3/287 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(132.71 30.52 132.84 30.67)
MU9413/3/reg_r_shiftReg_44_/1 G_DG U9413/3/CLK U9413/3/271 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(115.485 30.52 115.615 30.67)
MU9413/3/reg_r_shiftReg_44_/2 U9413/3/272 U9413/3/271 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(116.065 30.52 116.195 30.67)
MU9413/3/reg_r_shiftReg_44_/3 U9413/3/reg_r_shiftReg_44_/4 U9413/3/ix1816/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(117.155 30.52 117.285 30.67)
MU9413/3/reg_r_shiftReg_44_/4 U9413/3/275 U9413/3/271 U9413/3/reg_r_shiftReg_44_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(117.67 30.52 117.8 30.67)
MU9413/3/reg_r_shiftReg_44_/5 U9413/3/276 U9413/3/275 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(118.76 30.52 118.89 30.67)
MU9413/3/reg_r_shiftReg_44_/6 U9413/3/reg_r_shiftReg_44_/7 U9413/3/CLB U9413/3/275 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(120.13 30.52 120.26 30.67)
MU9413/3/reg_r_shiftReg_44_/7 U9413/3/reg_r_shiftReg_44_/8 U9413/3/276 U9413/3/reg_r_shiftReg_44_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(120.61 30.52 120.74 30.67)
MU9413/3/reg_r_shiftReg_44_/8 G_DG U9413/3/272 U9413/3/reg_r_shiftReg_44_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(121.09 30.52 121.22 30.67)
MU9413/3/reg_r_shiftReg_44_/9 U9413/3/reg_r_shiftReg_44_/9 U9413/3/276 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(122.18 30.52 122.31 30.67)
MU9413/3/reg_r_shiftReg_44_/10 U9413/3/reg_r_shiftReg_44_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_44_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(122.69 30.52 122.82 30.67)
MU9413/3/reg_r_shiftReg_44_/11 U9413/3/279 U9413/3/272 U9413/3/reg_r_shiftReg_44_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(123.11 30.52 123.24 30.67)
MU9413/3/reg_r_shiftReg_44_/12 U9413/3/280 U9413/3/279 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(124.2 30.52 124.33 30.67)
MU9413/3/reg_r_shiftReg_44_/13 U9413/3/281 U9413/3/271 U9413/3/279 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(125.56 30.52 125.69 30.67)
MU9413/3/reg_r_shiftReg_44_/14 U9413/3/reg_r_shiftReg_44_/14 U9413/3/CLB U9413/3/281 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(126.14 30.52 126.27 30.67)
MU9413/3/reg_r_shiftReg_44_/15 G_DG U9413/3/280 U9413/3/reg_r_shiftReg_44_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(126.45 30.52 126.58 30.67)
MU9413/3/reg_r_shiftReg_44_/16 addr[11] U9413/3/281 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(127.54 30.52 127.67 30.67)
MU9413/3/reg_r_shiftReg_44_/17 U9413/3/reg_r_shiftReg_44_/QB U9413/3/280 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(128.63 30.52 128.76 30.67)
MU9413/3/ix2187/1 U9413/3/ix2187/1 rdData[2] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(112.565 30.52 112.695 30.67)
MU9413/3/ix2187/2 U9413/3/ix2187/OUT U9413/2/ix1948/B U9413/3/ix2187/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(113.145 30.52 113.275 30.67)
MU9413/3/ix2187/3 U9413/3/ix2187/3 wrData[2] U9413/3/ix2187/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(113.725 30.52 113.855 30.67)
MU9413/3/ix2187/4 G_DG U9413/D U9413/3/ix2187/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(114.305 30.52 114.435 30.67)
MU9413/3/ix85/1 U9413/3/ix85/1 U9413/3/ix2187/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(110.805 30.52 110.935 30.67)
MU9413/3/ix85/2 U9413/ix1786\Cross U9413/2/ix2189/OUT U9413/3/ix85/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(111.385 30.52 111.515 30.67)
MU9413/3/ix2181/1 U9413/3/ix2181/1 rdData[3] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(107.885 30.52 108.015 30.67)
MU9413/3/ix2181/2 U9413/3/ix2181/OUT U9413/2/ix1948/B U9413/3/ix2181/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(108.465 30.52 108.595 30.67)
MU9413/3/ix2181/3 U9413/3/ix2181/3 wrData[3] U9413/3/ix2181/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(109.045 30.52 109.175 30.67)
MU9413/3/ix2181/4 G_DG U9413/D U9413/3/ix2181/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(109.625 30.52 109.755 30.67)
MU9413/3/ix2177/1 U9413/3/ix2177/1 wrData[3] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(106.125 30.52 106.255 30.67)
MU9413/3/ix2177/2 U9413/3/ix109/B U9413/2/ix2147/B U9413/3/ix2177/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(106.705 30.52 106.835 30.67)
MU9413/3/ix109/1 U9413/3/ix109/1 U9413/2/ix2175/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(104.365 30.52 104.495 30.67)
MU9413/3/ix109/2 U9413/3/ix109/OUT U9413/3/ix109/B U9413/3/ix109/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(104.945 30.52 105.075 30.67)
MU9413/3/reg_r_shiftReg_5_/1 G_DG U9413/3/CLK U9413/3/239 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(90.04 30.52 90.17 30.67)
MU9413/3/reg_r_shiftReg_5_/2 U9413/3/240 U9413/3/239 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(90.62 30.52 90.75 30.67)
MU9413/3/reg_r_shiftReg_5_/3 U9413/3/reg_r_shiftReg_5_/4 U9413/3/ix109/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(91.71 30.52 91.84 30.67)
MU9413/3/reg_r_shiftReg_5_/4 U9413/3/243 U9413/3/239 U9413/3/reg_r_shiftReg_5_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(92.225 30.52 92.355 30.67)
MU9413/3/reg_r_shiftReg_5_/5 U9413/3/244 U9413/3/243 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(93.315 30.52 93.445 30.67)
MU9413/3/reg_r_shiftReg_5_/6 U9413/3/reg_r_shiftReg_5_/7 U9413/3/CLB U9413/3/243 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(94.685 30.52 94.815 30.67)
MU9413/3/reg_r_shiftReg_5_/7 U9413/3/reg_r_shiftReg_5_/8 U9413/3/244 U9413/3/reg_r_shiftReg_5_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(95.165 30.52 95.295 30.67)
MU9413/3/reg_r_shiftReg_5_/8 G_DG U9413/3/240 U9413/3/reg_r_shiftReg_5_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(95.645 30.52 95.775 30.67)
MU9413/3/reg_r_shiftReg_5_/9 U9413/3/reg_r_shiftReg_5_/9 U9413/3/244 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(96.735 30.52 96.865 30.67)
MU9413/3/reg_r_shiftReg_5_/10 U9413/3/reg_r_shiftReg_5_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_5_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(97.245 30.52 97.375 30.67)
MU9413/3/reg_r_shiftReg_5_/11 U9413/3/247 U9413/3/240 U9413/3/reg_r_shiftReg_5_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(97.665 30.52 97.795 30.67)
MU9413/3/reg_r_shiftReg_5_/12 U9413/3/248 U9413/3/247 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(98.755 30.52 98.885 30.67)
MU9413/3/reg_r_shiftReg_5_/13 U9413/3/249 U9413/3/239 U9413/3/247 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(100.115 30.52 100.245 30.67)
MU9413/3/reg_r_shiftReg_5_/14 U9413/3/reg_r_shiftReg_5_/14 U9413/3/CLB U9413/3/249 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(100.695 30.52 100.825 30.67)
MU9413/3/reg_r_shiftReg_5_/15 G_DG U9413/3/248 U9413/3/reg_r_shiftReg_5_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(101.005 30.52 101.135 30.67)
MU9413/3/reg_r_shiftReg_5_/16 wrData[4] U9413/3/249 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(102.095 30.52 102.225 30.67)
MU9413/3/reg_r_shiftReg_5_/17 U9413/3/reg_r_shiftReg_5_/QB U9413/3/248 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(103.185 30.52 103.315 30.67)
MU9413/3/ix2165/1 U9413/3/ix2165/1 wrData[5] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(88.28 30.52 88.41 30.67)
MU9413/3/ix2165/2 U9413/3/ix133/B U9413/2/ix2147/B U9413/3/ix2165/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(88.86 30.52 88.99 30.67)
MU9413/3/ix2163/1 U9413/3/ix2163/1 rdData[6] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(85.36 30.52 85.49 30.67)
MU9413/3/ix2163/2 U9413/3/ix133/A U9413/2/ix2121/B U9413/3/ix2163/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(85.94 30.52 86.07 30.67)
MU9413/3/ix2163/3 U9413/3/ix2163/3 wrData[6] U9413/3/ix133/A G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(86.52 30.52 86.65 30.67)
MU9413/3/ix2163/4 G_DG U9413/2/ix2121/D U9413/3/ix2163/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(87.1 30.52 87.23 30.67)
MU9413/3/ix133/1 U9413/3/ix133/1 U9413/3/ix133/A G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(83.6 30.52 83.73 30.67)
MU9413/3/ix133/2 U9413/3/ix133/OUT U9413/3/ix133/B U9413/3/ix133/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(84.18 30.52 84.31 30.67)
MU9413/3/ix2296/1 G_DG U9413/3/ix2292/A U9413/3/225 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(81.84 30.52 81.97 30.67)
MU9413/3/ix2296/2 U9413/2/ix1948/B U9413/3/225 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(82.42 30.52 82.55 30.67)
MU9413/3/ix2157/1 U9413/3/ix2157/1 rdData[7] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(78.92 30.52 79.05 30.67)
MU9413/3/ix2157/2 U9413/3/ix2157/OUT U9413/2/ix2121/B U9413/3/ix2157/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(79.5 30.52 79.63 30.67)
MU9413/3/ix2157/3 U9413/3/ix2157/3 wrData[7] U9413/3/ix2157/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(80.08 30.52 80.21 30.67)
MU9413/3/ix2157/4 G_DG U9413/2/ix2121/D U9413/3/ix2157/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(80.66 30.52 80.79 30.67)
MU9413/3/ix2151/1 U9413/3/ix2151/1 rdData[8] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(76 30.52 76.13 30.67)
MU9413/3/ix2151/2 U9413/3/ix2151/OUT U9413/2/ix2121/B U9413/3/ix2151/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(76.58 30.52 76.71 30.67)
MU9413/3/ix2151/3 U9413/3/ix2151/3 wrData[8] U9413/3/ix2151/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(77.16 30.52 77.29 30.67)
MU9413/3/ix2151/4 G_DG U9413/2/ix2121/D U9413/3/ix2151/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(77.74 30.52 77.87 30.67)
MU9413/3/reg_r_shiftReg_11_/1 G_DG U9413/3/CLK U9413/3/199 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(61.675 30.52 61.805 30.67)
MU9413/3/reg_r_shiftReg_11_/2 U9413/3/200 U9413/3/199 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(62.255 30.52 62.385 30.67)
MU9413/3/reg_r_shiftReg_11_/3 U9413/3/reg_r_shiftReg_11_/4 U9413/2/ix181/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(63.345 30.52 63.475 30.67)
MU9413/3/reg_r_shiftReg_11_/4 U9413/3/203 U9413/3/199 U9413/3/reg_r_shiftReg_11_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(63.86 30.52 63.99 30.67)
MU9413/3/reg_r_shiftReg_11_/5 U9413/3/204 U9413/3/203 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(64.95 30.52 65.08 30.67)
MU9413/3/reg_r_shiftReg_11_/6 U9413/3/reg_r_shiftReg_11_/7 U9413/3/CLB U9413/3/203 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(66.32 30.52 66.45 30.67)
MU9413/3/reg_r_shiftReg_11_/7 U9413/3/reg_r_shiftReg_11_/8 U9413/3/204 U9413/3/reg_r_shiftReg_11_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(66.8 30.52 66.93 30.67)
MU9413/3/reg_r_shiftReg_11_/8 G_DG U9413/3/200 U9413/3/reg_r_shiftReg_11_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(67.28 30.52 67.41 30.67)
MU9413/3/reg_r_shiftReg_11_/9 U9413/3/reg_r_shiftReg_11_/9 U9413/3/204 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(68.37 30.52 68.5 30.67)
MU9413/3/reg_r_shiftReg_11_/10 U9413/3/reg_r_shiftReg_11_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_11_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(68.88 30.52 69.01 30.67)
MU9413/3/reg_r_shiftReg_11_/11 U9413/3/207 U9413/3/200 U9413/3/reg_r_shiftReg_11_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(69.3 30.52 69.43 30.67)
MU9413/3/reg_r_shiftReg_11_/12 U9413/3/208 U9413/3/207 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(70.39 30.52 70.52 30.67)
MU9413/3/reg_r_shiftReg_11_/13 U9413/3/209 U9413/3/199 U9413/3/207 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(71.75 30.52 71.88 30.67)
MU9413/3/reg_r_shiftReg_11_/14 U9413/3/reg_r_shiftReg_11_/14 U9413/3/CLB U9413/3/209 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(72.33 30.52 72.46 30.67)
MU9413/3/reg_r_shiftReg_11_/15 G_DG U9413/3/208 U9413/3/reg_r_shiftReg_11_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(72.64 30.52 72.77 30.67)
MU9413/3/reg_r_shiftReg_11_/16 wrData[10] U9413/3/209 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(73.73 30.52 73.86 30.67)
MU9413/3/reg_r_shiftReg_11_/17 U9413/3/reg_r_shiftReg_11_/QB U9413/3/208 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(74.82 30.52 74.95 30.67)
MU9413/3/ix2135/1 U9413/3/ix2135/1 wrData[10] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(59.915 30.52 60.045 30.67)
MU9413/3/ix2135/2 U9413/3/ix193/B U9413/2/ix2093/B U9413/3/ix2135/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(60.495 30.52 60.625 30.67)
MU9413/3/ix193/1 U9413/3/ix193/1 U9413/2/ix2133/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(58.155 30.52 58.285 30.67)
MU9413/3/ix193/2 U9413/3/ix193/OUT U9413/3/ix193/B U9413/3/ix193/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(58.735 30.52 58.865 30.67)
MU9413/3/ix2294/1 G_DG U9413/3/ix2292/A U9413/3/191 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(56.395 30.52 56.525 30.67)
MU9413/3/ix2294/2 U9413/2/ix2121/B U9413/3/191 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(56.975 30.52 57.105 30.67)
MU9413/3/ix2123/1 U9413/3/ix2123/1 wrData[12] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(54.635 30.52 54.765 30.67)
MU9413/3/ix2123/2 U9413/3/ix2123/OUT U9413/2/ix2093/B U9413/3/ix2123/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(55.215 30.52 55.345 30.67)
MU9413/3/ix217/1 U9413/3/ix217/1 U9413/2/ix2121/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(52.875 30.52 53.005 30.67)
MU9413/3/ix217/2 U9413/3/ix217/OUT U9413/3/ix2123/OUT U9413/3/ix217/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(53.455 30.52 53.585 30.67)
MU9413/3/reg_r_shiftReg_17_/1 G_DG U9413/3/CLK U9413/3/171 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(38.55 30.52 38.68 30.67)
MU9413/3/reg_r_shiftReg_17_/2 U9413/3/172 U9413/3/171 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(39.13 30.52 39.26 30.67)
MU9413/3/reg_r_shiftReg_17_/3 U9413/3/reg_r_shiftReg_17_/4 U9413/3/ix253/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(40.22 30.52 40.35 30.67)
MU9413/3/reg_r_shiftReg_17_/4 U9413/3/175 U9413/3/171 U9413/3/reg_r_shiftReg_17_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(40.735 30.52 40.865 30.67)
MU9413/3/reg_r_shiftReg_17_/5 U9413/3/176 U9413/3/175 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(41.825 30.52 41.955 30.67)
MU9413/3/reg_r_shiftReg_17_/6 U9413/3/reg_r_shiftReg_17_/7 U9413/3/CLB U9413/3/175 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(43.195 30.52 43.325 30.67)
MU9413/3/reg_r_shiftReg_17_/7 U9413/3/reg_r_shiftReg_17_/8 U9413/3/176 U9413/3/reg_r_shiftReg_17_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(43.675 30.52 43.805 30.67)
MU9413/3/reg_r_shiftReg_17_/8 G_DG U9413/3/172 U9413/3/reg_r_shiftReg_17_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(44.155 30.52 44.285 30.67)
MU9413/3/reg_r_shiftReg_17_/9 U9413/3/reg_r_shiftReg_17_/9 U9413/3/176 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(45.245 30.52 45.375 30.67)
MU9413/3/reg_r_shiftReg_17_/10 U9413/3/reg_r_shiftReg_17_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_17_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(45.755 30.52 45.885 30.67)
MU9413/3/reg_r_shiftReg_17_/11 U9413/3/179 U9413/3/172 U9413/3/reg_r_shiftReg_17_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(46.175 30.52 46.305 30.67)
MU9413/3/reg_r_shiftReg_17_/12 U9413/3/180 U9413/3/179 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(47.265 30.52 47.395 30.67)
MU9413/3/reg_r_shiftReg_17_/13 U9413/3/181 U9413/3/171 U9413/3/179 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(48.625 30.52 48.755 30.67)
MU9413/3/reg_r_shiftReg_17_/14 U9413/3/reg_r_shiftReg_17_/14 U9413/3/CLB U9413/3/181 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(49.205 30.52 49.335 30.67)
MU9413/3/reg_r_shiftReg_17_/15 G_DG U9413/3/180 U9413/3/reg_r_shiftReg_17_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(49.515 30.52 49.645 30.67)
MU9413/3/reg_r_shiftReg_17_/16 wrData[16] U9413/3/181 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(50.605 30.52 50.735 30.67)
MU9413/3/reg_r_shiftReg_17_/17 U9413/3/reg_r_shiftReg_17_/QB U9413/3/180 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(51.695 30.52 51.825 30.67)
MU9413/3/ix253/1 U9413/3/ix253/1 U9413/3/ix2103/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(36.79 30.52 36.92 30.67)
MU9413/3/ix253/2 U9413/3/ix253/OUT U9413/2/ix2105/OUT U9413/3/ix253/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(37.37 30.52 37.5 30.67)
MU9413/3/ix2115/1 U9413/3/ix2115/1 rdData[14] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(33.87 30.52 34 30.67)
MU9413/3/ix2115/2 U9413/3/ix2115/OUT U9413/2/ix2067/B U9413/3/ix2115/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(34.45 30.52 34.58 30.67)
MU9413/3/ix2115/3 U9413/3/ix2115/3 wrData[14] U9413/3/ix2115/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(35.03 30.52 35.16 30.67)
MU9413/3/ix2115/4 G_DG U9413/2/ix2067/D U9413/3/ix2115/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(35.61 30.52 35.74 30.67)
MU9413/3/ix2103/1 U9413/3/ix2103/1 rdData[16] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(30.95 30.52 31.08 30.67)
MU9413/3/ix2103/2 U9413/3/ix2103/OUT U9413/2/ix2067/B U9413/3/ix2103/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(31.53 30.52 31.66 30.67)
MU9413/3/ix2103/3 U9413/3/ix2103/3 wrData[16] U9413/3/ix2103/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(32.11 30.52 32.24 30.67)
MU9413/3/ix2103/4 G_DG U9413/2/ix2067/D U9413/3/ix2103/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(32.69 30.52 32.82 30.67)
MU9413/3/reg_r_shiftReg_20_/1 G_DG U9413/3/CLK U9413/3/143 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(16.625 30.52 16.755 30.67)
MU9413/3/reg_r_shiftReg_20_/2 U9413/3/144 U9413/3/143 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(17.205 30.52 17.335 30.67)
MU9413/3/reg_r_shiftReg_20_/3 U9413/3/reg_r_shiftReg_20_/4 U9413/2/ix289/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(18.295 30.52 18.425 30.67)
MU9413/3/reg_r_shiftReg_20_/4 U9413/3/147 U9413/3/143 U9413/3/reg_r_shiftReg_20_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(18.81 30.52 18.94 30.67)
MU9413/3/reg_r_shiftReg_20_/5 U9413/3/148 U9413/3/147 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(19.9 30.52 20.03 30.67)
MU9413/3/reg_r_shiftReg_20_/6 U9413/3/reg_r_shiftReg_20_/7 U9413/3/CLB U9413/3/147 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(21.27 30.52 21.4 30.67)
MU9413/3/reg_r_shiftReg_20_/7 U9413/3/reg_r_shiftReg_20_/8 U9413/3/148 U9413/3/reg_r_shiftReg_20_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(21.75 30.52 21.88 30.67)
MU9413/3/reg_r_shiftReg_20_/8 G_DG U9413/3/144 U9413/3/reg_r_shiftReg_20_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(22.23 30.52 22.36 30.67)
MU9413/3/reg_r_shiftReg_20_/9 U9413/3/reg_r_shiftReg_20_/9 U9413/3/148 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(23.32 30.52 23.45 30.67)
MU9413/3/reg_r_shiftReg_20_/10 U9413/3/reg_r_shiftReg_20_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_20_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(23.83 30.52 23.96 30.67)
MU9413/3/reg_r_shiftReg_20_/11 U9413/3/151 U9413/3/144 U9413/3/reg_r_shiftReg_20_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(24.25 30.52 24.38 30.67)
MU9413/3/reg_r_shiftReg_20_/12 U9413/3/152 U9413/3/151 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(25.34 30.52 25.47 30.67)
MU9413/3/reg_r_shiftReg_20_/13 U9413/3/153 U9413/3/143 U9413/3/151 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(26.7 30.52 26.83 30.67)
MU9413/3/reg_r_shiftReg_20_/14 U9413/3/reg_r_shiftReg_20_/14 U9413/3/CLB U9413/3/153 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(27.28 30.52 27.41 30.67)
MU9413/3/reg_r_shiftReg_20_/15 G_DG U9413/3/152 U9413/3/reg_r_shiftReg_20_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(27.59 30.52 27.72 30.67)
MU9413/3/reg_r_shiftReg_20_/16 wrData[19] U9413/3/153 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(28.68 30.52 28.81 30.67)
MU9413/3/reg_r_shiftReg_20_/17 U9413/3/reg_r_shiftReg_20_/QB U9413/3/152 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(29.77 30.52 29.9 30.67)
MU9413/3/ix2097/1 U9413/3/ix2097/1 rdData[17] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(13.705 30.52 13.835 30.67)
MU9413/3/ix2097/2 U9413/3/ix2097/OUT U9413/2/ix2067/B U9413/3/ix2097/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(14.285 30.52 14.415 30.67)
MU9413/3/ix2097/3 U9413/3/ix2097/3 wrData[17] U9413/3/ix2097/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(14.865 30.52 14.995 30.67)
MU9413/3/ix2097/4 G_DG U9413/2/ix2067/D U9413/3/ix2097/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(15.445 30.52 15.575 30.67)
MU9413/3/ix2292/1 G_DG U9413/3/ix2292/A U9413/3/135 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(11.945 30.52 12.075 30.67)
MU9413/3/ix2292/2 U9413/2/ix2067/B U9413/3/135 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(12.525 30.52 12.655 30.67)
MU9413/3/ix2081/1 U9413/3/ix2081/1 wrData[19] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(10.185 30.52 10.315 30.67)
MU9413/3/ix2081/2 U9413/3/ix2081/OUT U9413/2/ix2045/B U9413/3/ix2081/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(10.765 30.52 10.895 30.67)
MU9413/3/ix301/1 U9413/3/ix301/1 U9413/2/ix2079/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(8.425 30.52 8.555 30.67)
MU9413/3/ix301/2 U9413/3/ix301/OUT U9413/3/ix2081/OUT U9413/3/ix301/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(9.005 30.52 9.135 30.67)
MU9413/3/reg_r_shiftReg_21_/1 G_DG U9413/3/CLK U9413/3/115 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-5.9 30.52 -5.77 30.67)
MU9413/3/reg_r_shiftReg_21_/2 U9413/3/116 U9413/3/115 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-5.32 30.52 -5.19 30.67)
MU9413/3/reg_r_shiftReg_21_/3 U9413/3/reg_r_shiftReg_21_/4 U9413/3/ix301/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-4.23 30.52 -4.1 30.67)
MU9413/3/reg_r_shiftReg_21_/4 U9413/3/119 U9413/3/115 U9413/3/reg_r_shiftReg_21_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-3.715 30.52 -3.585 30.67)
MU9413/3/reg_r_shiftReg_21_/5 U9413/3/120 U9413/3/119 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-2.625 30.52 -2.495 30.67)
MU9413/3/reg_r_shiftReg_21_/6 U9413/3/reg_r_shiftReg_21_/7 U9413/3/CLB U9413/3/119 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-1.255 30.52 -1.125 30.67)
MU9413/3/reg_r_shiftReg_21_/7 U9413/3/reg_r_shiftReg_21_/8 U9413/3/120 U9413/3/reg_r_shiftReg_21_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-0.775 30.52 -0.645 30.67)
MU9413/3/reg_r_shiftReg_21_/8 G_DG U9413/3/116 U9413/3/reg_r_shiftReg_21_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-0.295 30.52 -0.165 30.67)
MU9413/3/reg_r_shiftReg_21_/9 U9413/3/reg_r_shiftReg_21_/9 U9413/3/120 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(0.795 30.52 0.925 30.67)
MU9413/3/reg_r_shiftReg_21_/10 U9413/3/reg_r_shiftReg_21_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_21_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(1.305 30.52 1.435 30.67)
MU9413/3/reg_r_shiftReg_21_/11 U9413/3/123 U9413/3/116 U9413/3/reg_r_shiftReg_21_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(1.725 30.52 1.855 30.67)
MU9413/3/reg_r_shiftReg_21_/12 U9413/3/124 U9413/3/123 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(2.815 30.52 2.945 30.67)
MU9413/3/reg_r_shiftReg_21_/13 U9413/3/125 U9413/3/115 U9413/3/123 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(4.175 30.52 4.305 30.67)
MU9413/3/reg_r_shiftReg_21_/14 U9413/3/reg_r_shiftReg_21_/14 U9413/3/CLB U9413/3/125 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(4.755 30.52 4.885 30.67)
MU9413/3/reg_r_shiftReg_21_/15 G_DG U9413/3/124 U9413/3/reg_r_shiftReg_21_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(5.065 30.52 5.195 30.67)
MU9413/3/reg_r_shiftReg_21_/16 wrData[20] U9413/3/125 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(6.155 30.52 6.285 30.67)
MU9413/3/reg_r_shiftReg_21_/17 U9413/3/reg_r_shiftReg_21_/QB U9413/3/124 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(7.245 30.52 7.375 30.67)
MU9413/3/ix2073/1 U9413/3/ix2073/1 rdData[21] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-8.82 30.52 -8.69 30.67)
MU9413/3/ix2073/2 U9413/3/ix2073/OUT U9413/2/ix2067/B U9413/3/ix2073/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-8.24 30.52 -8.11 30.67)
MU9413/3/ix2073/3 U9413/3/ix2073/3 wrData[21] U9413/3/ix2073/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-7.66 30.52 -7.53 30.67)
MU9413/3/ix2073/4 G_DG U9413/2/ix2067/D U9413/3/ix2073/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-7.08 30.52 -6.95 30.67)
MU9413/3/reg_r_shiftReg_24_/1 G_DG U9413/3/CLK U9413/3/96 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-23.145 30.52 -23.015 30.67)
MU9413/3/reg_r_shiftReg_24_/2 U9413/3/97 U9413/3/96 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-22.565 30.52 -22.435 30.67)
MU9413/3/reg_r_shiftReg_24_/3 U9413/3/reg_r_shiftReg_24_/4 U9413/3/ix337/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-21.475 30.52 -21.345 30.67)
MU9413/3/reg_r_shiftReg_24_/4 U9413/3/100 U9413/3/96 U9413/3/reg_r_shiftReg_24_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-20.96 30.52 -20.83 30.67)
MU9413/3/reg_r_shiftReg_24_/5 U9413/3/101 U9413/3/100 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-19.87 30.52 -19.74 30.67)
MU9413/3/reg_r_shiftReg_24_/6 U9413/3/reg_r_shiftReg_24_/7 U9413/3/CLB U9413/3/100 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-18.5 30.52 -18.37 30.67)
MU9413/3/reg_r_shiftReg_24_/7 U9413/3/reg_r_shiftReg_24_/8 U9413/3/101 U9413/3/reg_r_shiftReg_24_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-18.02 30.52 -17.89 30.67)
MU9413/3/reg_r_shiftReg_24_/8 G_DG U9413/3/97 U9413/3/reg_r_shiftReg_24_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-17.54 30.52 -17.41 30.67)
MU9413/3/reg_r_shiftReg_24_/9 U9413/3/reg_r_shiftReg_24_/9 U9413/3/101 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-16.45 30.52 -16.32 30.67)
MU9413/3/reg_r_shiftReg_24_/10 U9413/3/reg_r_shiftReg_24_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_24_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-15.94 30.52 -15.81 30.67)
MU9413/3/reg_r_shiftReg_24_/11 U9413/3/104 U9413/3/97 U9413/3/reg_r_shiftReg_24_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-15.52 30.52 -15.39 30.67)
MU9413/3/reg_r_shiftReg_24_/12 U9413/3/105 U9413/3/104 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-14.43 30.52 -14.3 30.67)
MU9413/3/reg_r_shiftReg_24_/13 U9413/3/106 U9413/3/96 U9413/3/104 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-13.07 30.52 -12.94 30.67)
MU9413/3/reg_r_shiftReg_24_/14 U9413/3/reg_r_shiftReg_24_/14 U9413/3/CLB U9413/3/106 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-12.49 30.52 -12.36 30.67)
MU9413/3/reg_r_shiftReg_24_/15 G_DG U9413/3/105 U9413/3/reg_r_shiftReg_24_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-12.18 30.52 -12.05 30.67)
MU9413/3/reg_r_shiftReg_24_/16 wrData[23] U9413/3/106 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-11.09 30.52 -10.96 30.67)
MU9413/3/reg_r_shiftReg_24_/17 U9413/3/reg_r_shiftReg_24_/QB U9413/3/105 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-10 30.52 -9.87 30.67)
MU9413/3/ix337/1 U9413/3/ix337/1 U9413/2/ix2061/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-24.905 30.52 -24.775 30.67)
MU9413/3/ix337/2 U9413/3/ix337/OUT U9413/3/ix2063/OUT U9413/3/ix337/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-24.325 30.52 -24.195 30.67)
MU9413/3/ix2063/1 U9413/3/ix2063/1 wrData[22] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-26.665 30.52 -26.535 30.67)
MU9413/3/ix2063/2 U9413/3/ix2063/OUT U9413/2/ix2045/B U9413/3/ix2063/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-26.085 30.52 -25.955 30.67)
MU9413/3/ix2057/1 U9413/3/ix2057/1 wrData[23] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-28.425 30.52 -28.295 30.67)
MU9413/3/ix2057/2 U9413/3/ix2057/OUT U9413/2/ix2045/B U9413/3/ix2057/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-27.845 30.52 -27.715 30.67)
MU9413/3/ix349/1 U9413/3/ix349/1 U9413/3/ix2055/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-30.185 30.52 -30.055 30.67)
MU9413/3/ix349/2 U9413/3/ix349/OUT U9413/3/ix2057/OUT U9413/3/ix349/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-29.605 30.52 -29.475 30.67)
MU9413/3/ix2055/1 U9413/3/ix2055/1 rdData[24] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-33.105 30.52 -32.975 30.67)
MU9413/3/ix2055/2 U9413/3/ix2055/OUT U9413/2/ix2019/B U9413/3/ix2055/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-32.525 30.52 -32.395 30.67)
MU9413/3/ix2055/3 U9413/3/ix2055/3 wrData[24] U9413/3/ix2055/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-31.945 30.52 -31.815 30.67)
MU9413/3/ix2055/4 G_DG U9413/2/ix2019/D U9413/3/ix2055/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-31.365 30.52 -31.235 30.67)
MU9413/3/reg_r_shiftReg_27_/1 G_DG U9413/3/CLK U9413/3/65 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-47.43 30.52 -47.3 30.67)
MU9413/3/reg_r_shiftReg_27_/2 U9413/3/66 U9413/3/65 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-46.85 30.52 -46.72 30.67)
MU9413/3/reg_r_shiftReg_27_/3 U9413/3/reg_r_shiftReg_27_/4 U9413/2/ix373/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-45.76 30.52 -45.63 30.67)
MU9413/3/reg_r_shiftReg_27_/4 U9413/3/69 U9413/3/65 U9413/3/reg_r_shiftReg_27_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-45.245 30.52 -45.115 30.67)
MU9413/3/reg_r_shiftReg_27_/5 U9413/3/70 U9413/3/69 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-44.155 30.52 -44.025 30.67)
MU9413/3/reg_r_shiftReg_27_/6 U9413/3/reg_r_shiftReg_27_/7 U9413/3/CLB U9413/3/69 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-42.785 30.52 -42.655 30.67)
MU9413/3/reg_r_shiftReg_27_/7 U9413/3/reg_r_shiftReg_27_/8 U9413/3/70 U9413/3/reg_r_shiftReg_27_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-42.305 30.52 -42.175 30.67)
MU9413/3/reg_r_shiftReg_27_/8 G_DG U9413/3/66 U9413/3/reg_r_shiftReg_27_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-41.825 30.52 -41.695 30.67)
MU9413/3/reg_r_shiftReg_27_/9 U9413/3/reg_r_shiftReg_27_/9 U9413/3/70 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-40.735 30.52 -40.605 30.67)
MU9413/3/reg_r_shiftReg_27_/10 U9413/3/reg_r_shiftReg_27_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_27_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-40.225 30.52 -40.095 30.67)
MU9413/3/reg_r_shiftReg_27_/11 U9413/3/73 U9413/3/66 U9413/3/reg_r_shiftReg_27_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-39.805 30.52 -39.675 30.67)
MU9413/3/reg_r_shiftReg_27_/12 U9413/3/74 U9413/3/73 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-38.715 30.52 -38.585 30.67)
MU9413/3/reg_r_shiftReg_27_/13 U9413/3/75 U9413/3/65 U9413/3/73 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-37.355 30.52 -37.225 30.67)
MU9413/3/reg_r_shiftReg_27_/14 U9413/3/reg_r_shiftReg_27_/14 U9413/3/CLB U9413/3/75 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-36.775 30.52 -36.645 30.67)
MU9413/3/reg_r_shiftReg_27_/15 G_DG U9413/3/74 U9413/3/reg_r_shiftReg_27_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-36.465 30.52 -36.335 30.67)
MU9413/3/reg_r_shiftReg_27_/16 wrData[26] U9413/3/75 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-35.375 30.52 -35.245 30.67)
MU9413/3/reg_r_shiftReg_27_/17 U9413/3/reg_r_shiftReg_27_/QB U9413/3/74 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-34.285 30.52 -34.155 30.67)
MU9413/3/ix2039/1 U9413/3/ix2039/1 wrData[26] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-49.19 30.52 -49.06 30.67)
MU9413/3/ix2039/2 U9413/3/ix2039/OUT U9413/2/ix2045/B U9413/3/ix2039/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-48.61 30.52 -48.48 30.67)
MU9413/3/ix385/1 U9413/3/ix385/1 U9413/3/ix2037/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-50.95 30.52 -50.82 30.67)
MU9413/3/ix385/2 U9413/3/ix385/OUT U9413/3/ix2039/OUT U9413/3/ix385/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-50.37 30.52 -50.24 30.67)
MU9413/3/ix2037/1 U9413/3/ix2037/1 rdData[27] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-53.87 30.52 -53.74 30.67)
MU9413/3/ix2037/2 U9413/3/ix2037/OUT U9413/2/ix2019/B U9413/3/ix2037/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-53.29 30.52 -53.16 30.67)
MU9413/3/ix2037/3 U9413/3/ix2037/3 wrData[27] U9413/3/ix2037/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-52.71 30.52 -52.58 30.67)
MU9413/3/ix2037/4 G_DG U9413/2/ix2019/D U9413/3/ix2037/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-52.13 30.52 -52 30.67)
MU9413/3/reg_r_shiftReg_32_/1 G_DG U9413/3/CLK U9413/3/40 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-68.195 30.52 -68.065 30.67)
MU9413/3/reg_r_shiftReg_32_/2 U9413/3/41 U9413/3/40 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-67.615 30.52 -67.485 30.67)
MU9413/3/reg_r_shiftReg_32_/3 U9413/3/reg_r_shiftReg_32_/4 U9413/3/ix433/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-66.525 30.52 -66.395 30.67)
MU9413/3/reg_r_shiftReg_32_/4 U9413/3/44 U9413/3/40 U9413/3/reg_r_shiftReg_32_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-66.01 30.52 -65.88 30.67)
MU9413/3/reg_r_shiftReg_32_/5 U9413/3/45 U9413/3/44 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-64.92 30.52 -64.79 30.67)
MU9413/3/reg_r_shiftReg_32_/6 U9413/3/reg_r_shiftReg_32_/7 U9413/3/CLB U9413/3/44 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-63.55 30.52 -63.42 30.67)
MU9413/3/reg_r_shiftReg_32_/7 U9413/3/reg_r_shiftReg_32_/8 U9413/3/45 U9413/3/reg_r_shiftReg_32_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-63.07 30.52 -62.94 30.67)
MU9413/3/reg_r_shiftReg_32_/8 G_DG U9413/3/41 U9413/3/reg_r_shiftReg_32_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-62.59 30.52 -62.46 30.67)
MU9413/3/reg_r_shiftReg_32_/9 U9413/3/reg_r_shiftReg_32_/9 U9413/3/45 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-61.5 30.52 -61.37 30.67)
MU9413/3/reg_r_shiftReg_32_/10 U9413/3/reg_r_shiftReg_32_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_32_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-60.99 30.52 -60.86 30.67)
MU9413/3/reg_r_shiftReg_32_/11 U9413/3/48 U9413/3/41 U9413/3/reg_r_shiftReg_32_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-60.57 30.52 -60.44 30.67)
MU9413/3/reg_r_shiftReg_32_/12 U9413/3/49 U9413/3/48 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-59.48 30.52 -59.35 30.67)
MU9413/3/reg_r_shiftReg_32_/13 U9413/3/50 U9413/3/40 U9413/3/48 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-58.12 30.52 -57.99 30.67)
MU9413/3/reg_r_shiftReg_32_/14 U9413/3/reg_r_shiftReg_32_/14 U9413/3/CLB U9413/3/50 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-57.54 30.52 -57.41 30.67)
MU9413/3/reg_r_shiftReg_32_/15 G_DG U9413/3/49 U9413/3/reg_r_shiftReg_32_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-57.23 30.52 -57.1 30.67)
MU9413/3/reg_r_shiftReg_32_/16 wrData[31] U9413/3/50 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-56.14 30.52 -56.01 30.67)
MU9413/3/reg_r_shiftReg_32_/17 U9413/3/reg_r_shiftReg_32_/QB U9413/3/49 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-55.05 30.52 -54.92 30.67)
MU9413/3/ix2027/1 U9413/3/ix2027/1 wrData[28] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-69.955 30.52 -69.825 30.67)
MU9413/3/ix2027/2 U9413/3/ix2027/OUT U9413/2/ix2021/B U9413/3/ix2027/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-69.375 30.52 -69.245 30.67)
MU9413/3/ix433/1 U9413/3/ix433/1 U9413/3/ix1993/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-71.715 30.52 -71.585 30.67)
MU9413/3/ix433/2 U9413/3/ix433/OUT U9413/3/ix2015/OUT U9413/3/ix433/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-71.135 30.52 -71.005 30.67)
MU9413/3/ix2015/1 U9413/3/ix2015/1 wrData[30] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-73.475 30.52 -73.345 30.67)
MU9413/3/ix2015/2 U9413/3/ix2015/OUT U9413/2/ix2021/B U9413/3/ix2015/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-72.895 30.52 -72.765 30.67)
MU9413/3/ix1993/1 U9413/3/ix1993/1 rdData[31] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-76.395 30.52 -76.265 30.67)
MU9413/3/ix1993/2 U9413/3/ix1993/OUT U9413/2/ix2019/B U9413/3/ix1993/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-75.815 30.52 -75.685 30.67)
MU9413/3/ix1993/3 U9413/3/ix1993/3 wrData[31] U9413/3/ix1993/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-75.235 30.52 -75.105 30.67)
MU9413/3/ix1993/4 G_DG U9413/2/ix2019/D U9413/3/ix1993/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-74.655 30.52 -74.525 30.67)
MU9413/3/reg_r_shiftReg_47_/1 G_DG U9413/3/CLK U9413/3/12 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-90.72 30.52 -90.59 30.67)
MU9413/3/reg_r_shiftReg_47_/2 U9413/3/13 U9413/3/12 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-90.14 30.52 -90.01 30.67)
MU9413/3/reg_r_shiftReg_47_/3 U9413/3/reg_r_shiftReg_47_/4 U9413/3/ix1846/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-89.05 30.52 -88.92 30.67)
MU9413/3/reg_r_shiftReg_47_/4 U9413/3/16 U9413/3/12 U9413/3/reg_r_shiftReg_47_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-88.535 30.52 -88.405 30.67)
MU9413/3/reg_r_shiftReg_47_/5 U9413/3/17 U9413/3/16 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-87.445 30.52 -87.315 30.67)
MU9413/3/reg_r_shiftReg_47_/6 U9413/3/reg_r_shiftReg_47_/7 U9413/3/CLB U9413/3/16 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-86.075 30.52 -85.945 30.67)
MU9413/3/reg_r_shiftReg_47_/7 U9413/3/reg_r_shiftReg_47_/8 U9413/3/17 U9413/3/reg_r_shiftReg_47_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-85.595 30.52 -85.465 30.67)
MU9413/3/reg_r_shiftReg_47_/8 G_DG U9413/3/13 U9413/3/reg_r_shiftReg_47_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-85.115 30.52 -84.985 30.67)
MU9413/3/reg_r_shiftReg_47_/9 U9413/3/reg_r_shiftReg_47_/9 U9413/3/17 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-84.025 30.52 -83.895 30.67)
MU9413/3/reg_r_shiftReg_47_/10 U9413/3/reg_r_shiftReg_47_/10 U9413/3/CLB U9413/3/reg_r_shiftReg_47_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-83.515 30.52 -83.385 30.67)
MU9413/3/reg_r_shiftReg_47_/11 U9413/3/20 U9413/3/13 U9413/3/reg_r_shiftReg_47_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-83.095 30.52 -82.965 30.67)
MU9413/3/reg_r_shiftReg_47_/12 U9413/3/21 U9413/3/20 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-82.005 30.52 -81.875 30.67)
MU9413/3/reg_r_shiftReg_47_/13 U9413/3/22 U9413/3/12 U9413/3/20 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-80.645 30.52 -80.515 30.67)
MU9413/3/reg_r_shiftReg_47_/14 U9413/3/reg_r_shiftReg_47_/14 U9413/3/CLB U9413/3/22 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-80.065 30.52 -79.935 30.67)
MU9413/3/reg_r_shiftReg_47_/15 G_DG U9413/3/21 U9413/3/reg_r_shiftReg_47_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-79.755 30.52 -79.625 30.67)
MU9413/3/reg_r_shiftReg_47_/16 cmd[2] U9413/3/22 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-78.665 30.52 -78.535 30.67)
MU9413/3/reg_r_shiftReg_47_/17 U9413/3/reg_r_shiftReg_47_/QB U9413/3/21 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-77.575 30.52 -77.445 30.67)
MU9413/3/ix1846/1 G_DG U9413/SEL U9413/3/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-94.8 30.52 -94.67 30.67)
MU9413/3/ix1846/2 U9413/3/ix1846/3 U9413/3/5 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-94.22 30.52 -94.09 30.67)
MU9413/3/ix1846/3 U9413/3/7 cmd[2] U9413/3/ix1846/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-93.64 30.52 -93.51 30.67)
MU9413/3/ix1846/4 U9413/3/ix1846/5 cmd[1] U9413/3/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-93.06 30.52 -92.93 30.67)
MU9413/3/ix1846/5 G_DG U9413/SEL U9413/3/ix1846/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-92.48 30.52 -92.35 30.67)
MU9413/3/ix1846/6 U9413/3/ix1846/OUT U9413/3/7 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-91.9 30.52 -91.77 30.67)
MU9413/4/1 G_DS CLK U9413/4/2 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-98.32 21.715 -98.19 22.015)
MU9413/4/2 U9413/4/CLK U9413/4/2 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-97.74 21.715 -97.61 22.015)
MU9413/4/3 G_DS CLK U9413/4/3 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-96.56 21.715 -96.43 22.015)
MU9413/4/4 U9413/4/CLK U9413/4/3 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-95.98 21.715 -95.85 22.015)
MU9413/4/5 G_DS U9413/SEL U9413/4/5 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-94.8 21.5 -94.67 21.8)
MU9413/4/6 U9413/4/6 U9413/4/5 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-94.22 21.5 -94.09 22.02)
MU9413/4/7 U9413/4/7 cmd[0] U9413/4/6 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-93.64 21.5 -93.51 22.02)
MU9413/4/8 U9413/4/9 cmd[1] U9413/4/7 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-93.06 21.5 -92.93 22.02)
MU9413/4/9 G_DS U9413/SEL U9413/4/9 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-92.48 21.5 -92.35 22.02)
MU9413/4/10 U9413/4/ix1836/OUT U9413/4/7 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-91.9 21.715 -91.77 22.015)
MU9413/4/11 G_DS U9413/4/CLK U9413/4/12 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-90.72 21.715 -90.59 22.015)
MU9413/4/12 U9413/4/13 U9413/4/12 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-90.14 21.715 -90.01 22.015)
MU9413/4/13 U9413/4/14 U9413/4/ix1836/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-89.05 21.715 -88.92 22.105)
MU9413/4/14 U9413/4/16 U9413/4/13 U9413/4/14 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-88.535 21.715 -88.405 22.105)
MU9413/4/15 U9413/4/17 U9413/4/16 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-87.445 21.715 -87.315 22.015)
MU9413/4/16 U9413/4/18 U9413/4/12 U9413/4/16 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-86.355 21.715 -86.225 22.105)
MU9413/4/17 G_DS U9413/4/CLB U9413/4/18 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-85.735 21.715 -85.605 22.105)
MU9413/4/18 U9413/4/18 U9413/4/17 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-85.115 21.715 -84.985 22.105)
MU9413/4/19 U9413/4/19 U9413/4/17 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-84.025 21.715 -83.895 22.105)
MU9413/4/20 U9413/4/20 U9413/4/12 U9413/4/19 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-83.715 21.715 -83.585 22.105)
MU9413/4/21 U9413/4/21 U9413/4/20 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-82.005 21.715 -81.875 22.015)
MU9413/4/22 U9413/4/22 U9413/4/13 U9413/4/20 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-80.915 21.715 -80.785 22.105)
MU9413/4/23 G_DS U9413/4/CLB U9413/4/22 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-80.335 21.715 -80.205 22.105)
MU9413/4/24 U9413/4/22 U9413/4/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-79.755 21.715 -79.625 22.015)
MU9413/4/25 cmd[1] U9413/4/22 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-78.665 21.715 -78.535 22.015)
MU9413/4/26 U9413/4/reg_r_shiftReg_46_/QB U9413/4/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-77.575 21.715 -77.445 22.015)
MU9413/4/27 U9413/4/ix409/OUT U9413/reg_r_shiftReg_47_\Cross G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-76.395 21.715 -76.265 21.975)
MU9413/4/28 G_DS U9413/3/ix2027/OUT U9413/4/ix409/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-75.815 21.715 -75.685 21.975)
MU9413/4/29 G_DS U9413/4/CLK U9413/4/28 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-74.635 21.715 -74.505 22.015)
MU9413/4/30 U9413/4/29 U9413/4/28 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-74.055 21.715 -73.925 22.015)
MU9413/4/31 U9413/4/30 U9413/4/ix409/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-72.965 21.715 -72.835 22.105)
MU9413/4/32 U9413/4/32 U9413/4/29 U9413/4/30 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-72.45 21.715 -72.32 22.105)
MU9413/4/33 U9413/4/33 U9413/4/32 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-71.36 21.715 -71.23 22.015)
MU9413/4/34 U9413/4/34 U9413/4/28 U9413/4/32 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-70.27 21.715 -70.14 22.105)
MU9413/4/35 G_DS U9413/4/CLB U9413/4/34 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-69.65 21.715 -69.52 22.105)
MU9413/4/36 U9413/4/34 U9413/4/33 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-69.03 21.715 -68.9 22.105)
MU9413/4/37 U9413/4/35 U9413/4/33 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-67.94 21.715 -67.81 22.105)
MU9413/4/38 U9413/4/36 U9413/4/28 U9413/4/35 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-67.63 21.715 -67.5 22.105)
MU9413/4/39 U9413/4/37 U9413/4/36 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-65.92 21.715 -65.79 22.015)
MU9413/4/40 U9413/4/38 U9413/4/29 U9413/4/36 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-64.83 21.715 -64.7 22.105)
MU9413/4/41 G_DS U9413/4/CLB U9413/4/38 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-64.25 21.715 -64.12 22.105)
MU9413/4/42 U9413/4/38 U9413/4/37 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-63.67 21.715 -63.54 22.015)
MU9413/4/43 wrData[29] U9413/4/38 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-62.58 21.715 -62.45 22.015)
MU9413/4/44 U9413/4/reg_r_shiftReg_30_/QB U9413/4/37 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-61.49 21.715 -61.36 22.015)
MU9413/4/45 G_DS U9413/4/CLK U9413/4/41 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-60.31 21.715 -60.18 22.015)
MU9413/4/46 U9413/4/42 U9413/4/41 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-59.73 21.715 -59.6 22.015)
MU9413/4/47 U9413/4/43 U9413/3/ix385/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-58.64 21.715 -58.51 22.105)
MU9413/4/48 U9413/4/45 U9413/4/42 U9413/4/43 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-58.125 21.715 -57.995 22.105)
MU9413/4/49 U9413/4/46 U9413/4/45 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-57.035 21.715 -56.905 22.015)
MU9413/4/50 U9413/4/47 U9413/4/41 U9413/4/45 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-55.945 21.715 -55.815 22.105)
MU9413/4/51 G_DS U9413/4/CLB U9413/4/47 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-55.325 21.715 -55.195 22.105)
MU9413/4/52 U9413/4/47 U9413/4/46 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-54.705 21.715 -54.575 22.105)
MU9413/4/53 U9413/4/48 U9413/4/46 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-53.615 21.715 -53.485 22.105)
MU9413/4/54 U9413/4/49 U9413/4/41 U9413/4/48 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-53.305 21.715 -53.175 22.105)
MU9413/4/55 U9413/4/50 U9413/4/49 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-51.595 21.715 -51.465 22.015)
MU9413/4/56 U9413/4/51 U9413/4/42 U9413/4/49 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-50.505 21.715 -50.375 22.105)
MU9413/4/57 G_DS U9413/4/CLB U9413/4/51 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-49.925 21.715 -49.795 22.105)
MU9413/4/58 U9413/4/51 U9413/4/50 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-49.345 21.715 -49.215 22.015)
MU9413/4/59 wrData[27] U9413/4/51 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-48.255 21.715 -48.125 22.015)
MU9413/4/60 U9413/4/reg_r_shiftReg_28_/QB U9413/4/50 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-47.165 21.715 -47.035 22.015)
MU9413/4/61 G_DS U9413/4/CLK U9413/4/54 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-45.985 21.715 -45.855 22.015)
MU9413/4/62 U9413/4/55 U9413/4/54 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-45.405 21.715 -45.275 22.015)
MU9413/4/63 U9413/4/56 U9413/3/ix349/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-44.315 21.715 -44.185 22.105)
MU9413/4/64 U9413/4/58 U9413/4/55 U9413/4/56 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-43.8 21.715 -43.67 22.105)
MU9413/4/65 U9413/4/59 U9413/4/58 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-42.71 21.715 -42.58 22.015)
MU9413/4/66 U9413/4/60 U9413/4/54 U9413/4/58 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-41.62 21.715 -41.49 22.105)
MU9413/4/67 G_DS U9413/4/CLB U9413/4/60 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-41 21.715 -40.87 22.105)
MU9413/4/68 U9413/4/60 U9413/4/59 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-40.38 21.715 -40.25 22.105)
MU9413/4/69 U9413/4/61 U9413/4/59 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-39.29 21.715 -39.16 22.105)
MU9413/4/70 U9413/4/62 U9413/4/54 U9413/4/61 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-38.98 21.715 -38.85 22.105)
MU9413/4/71 U9413/4/63 U9413/4/62 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-37.27 21.715 -37.14 22.015)
MU9413/4/72 U9413/4/64 U9413/4/55 U9413/4/62 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-36.18 21.715 -36.05 22.105)
MU9413/4/73 G_DS U9413/4/CLB U9413/4/64 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-35.6 21.715 -35.47 22.105)
MU9413/4/74 U9413/4/64 U9413/4/63 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-35.02 21.715 -34.89 22.015)
MU9413/4/75 wrData[24] U9413/4/64 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-33.93 21.715 -33.8 22.015)
MU9413/4/76 U9413/4/reg_r_shiftReg_25_/QB U9413/4/63 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-32.84 21.715 -32.71 22.015)
MU9413/4/77 U9413/4/67 ack G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-31.66 21.5 -31.53 22.02)
MU9413/4/78 U9413/2/ix2019/D U9413/4/ix2270/OUT U9413/4/67 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-31.08 21.5 -30.95 22.02)
MU9413/4/79 G_DS U9413/4/ix2270/A U9413/4/72 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-29.9 21.715 -29.77 22.015)
MU9413/4/80 U9413/4/ix2270/OUT U9413/4/72 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-29.32 21.715 -29.19 22.015)
MU9413/4/81 G_DS U9413/4/CLK U9413/4/74 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-28.14 21.715 -28.01 22.015)
MU9413/4/82 U9413/4/75 U9413/4/74 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-27.56 21.715 -27.43 22.015)
MU9413/4/83 U9413/4/76 U9413/4/ix313/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-26.47 21.715 -26.34 22.105)
MU9413/4/84 U9413/4/78 U9413/4/75 U9413/4/76 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-25.955 21.715 -25.825 22.105)
MU9413/4/85 U9413/4/79 U9413/4/78 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-24.865 21.715 -24.735 22.015)
MU9413/4/86 U9413/4/80 U9413/4/74 U9413/4/78 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-23.775 21.715 -23.645 22.105)
MU9413/4/87 G_DS U9413/4/CLB U9413/4/80 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-23.155 21.715 -23.025 22.105)
MU9413/4/88 U9413/4/80 U9413/4/79 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-22.535 21.715 -22.405 22.105)
MU9413/4/89 U9413/4/81 U9413/4/79 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-21.445 21.715 -21.315 22.105)
MU9413/4/90 U9413/4/82 U9413/4/74 U9413/4/81 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-21.135 21.715 -21.005 22.105)
MU9413/4/91 U9413/4/83 U9413/4/82 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-19.425 21.715 -19.295 22.015)
MU9413/4/92 U9413/4/84 U9413/4/75 U9413/4/82 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-18.335 21.715 -18.205 22.105)
MU9413/4/93 G_DS U9413/4/CLB U9413/4/84 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-17.755 21.715 -17.625 22.105)
MU9413/4/94 U9413/4/84 U9413/4/83 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-17.175 21.715 -17.045 22.015)
MU9413/4/95 wrData[21] U9413/4/84 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-16.085 21.715 -15.955 22.015)
MU9413/4/96 U9413/4/reg_r_shiftReg_22_/QB U9413/4/83 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-14.995 21.715 -14.865 22.015)
MU9413/4/97 G_DS U9413/3/ix2292/A U9413/4/88 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-13.815 21.715 -13.685 22.015)
MU9413/4/98 U9413/2/ix2019/B U9413/4/88 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-13.235 21.715 -13.105 22.015)
MU9413/4/99 U9413/4/ix313/OUT U9413/3/ix2073/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-12.055 21.715 -11.925 21.975)
MU9413/4/100 G_DS U9413/4/ix2075/OUT U9413/4/ix313/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-11.475 21.715 -11.345 21.975)
MU9413/4/101 U9413/4/ix2075/OUT wrData[20] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-10.295 21.715 -10.165 21.975)
MU9413/4/102 G_DS U9413/2/ix2045/B U9413/4/ix2075/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-9.715 21.715 -9.585 21.975)
MU9413/4/103 U9413/4/96 ack G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-8.535 21.5 -8.405 22.02)
MU9413/4/104 U9413/2/ix2067/D U9413/4/ix2270/OUT U9413/4/96 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-7.955 21.5 -7.825 22.02)
MU9413/4/105 U9413/4/100 ack G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-6.775 21.5 -6.645 22.02)
MU9413/4/106 U9413/2/ix2121/D U9413/4/ix2270/OUT U9413/4/100 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-6.195 21.5 -6.065 22.02)
MU9413/4/107 G_DS U9413/4/ix2276/A U9413/4/105 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-5.015 21.715 -4.885 22.015)
MU9413/4/108 U9413/2/ix2021/B U9413/4/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-4.435 21.715 -4.305 22.015)
MU9413/4/109 G_DS U9413/4/ix2276/A U9413/4/108 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-3.255 21.715 -3.125 22.015)
MU9413/4/110 U9413/2/ix2045/B U9413/4/108 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-2.675 21.715 -2.545 22.015)
MU9413/4/111 U9413/reg_r_shiftReg_21_\Cross U9413/4/ix2251/A G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-1.495 21.715 -1.365 21.975)
MU9413/4/112 G_DS U9413/2/ix2021/B U9413/reg_r_shiftReg_21_\Cross G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-0.915 21.715 -0.785 21.975)
MU9413/4/113 G_DS U9413/4/CLK U9413/4/113 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(0.265 21.715 0.395 22.015)
MU9413/4/114 U9413/4/114 U9413/4/113 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(0.845 21.715 0.975 22.015)
MU9413/4/115 U9413/4/115 U9413/4/ix265/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(1.935 21.715 2.065 22.105)
MU9413/4/116 U9413/4/117 U9413/4/114 U9413/4/115 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(2.45 21.715 2.58 22.105)
MU9413/4/117 U9413/4/118 U9413/4/117 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(3.54 21.715 3.67 22.015)
MU9413/4/118 U9413/4/119 U9413/4/113 U9413/4/117 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(4.63 21.715 4.76 22.105)
MU9413/4/119 G_DS U9413/4/CLB U9413/4/119 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(5.25 21.715 5.38 22.105)
MU9413/4/120 U9413/4/119 U9413/4/118 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(5.87 21.715 6 22.105)
MU9413/4/121 U9413/4/120 U9413/4/118 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(6.96 21.715 7.09 22.105)
MU9413/4/122 U9413/4/121 U9413/4/113 U9413/4/120 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(7.27 21.715 7.4 22.105)
MU9413/4/123 U9413/4/122 U9413/4/121 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(8.98 21.715 9.11 22.015)
MU9413/4/124 U9413/4/123 U9413/4/114 U9413/4/121 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(10.07 21.715 10.2 22.105)
MU9413/4/125 G_DS U9413/4/CLB U9413/4/123 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(10.65 21.715 10.78 22.105)
MU9413/4/126 U9413/4/123 U9413/4/122 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(11.23 21.715 11.36 22.015)
MU9413/4/127 wrData[17] U9413/4/123 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(12.32 21.715 12.45 22.015)
MU9413/4/128 U9413/4/reg_r_shiftReg_18_/QB U9413/4/122 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(13.41 21.715 13.54 22.015)
MU9413/4/129 U9413/4/ix265/OUT U9413/3/ix2097/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(14.59 21.715 14.72 21.975)
MU9413/4/130 G_DS U9413/4/ix2099/OUT U9413/4/ix265/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(15.17 21.715 15.3 21.975)
MU9413/4/131 G_DS U9413/4/ix2276/A U9413/4/130 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(16.35 21.715 16.48 22.015)
MU9413/4/132 U9413/2/ix2093/B U9413/4/130 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(16.93 21.715 17.06 22.015)
MU9413/4/133 U9413/4/ix2099/OUT wrData[16] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(18.11 21.715 18.24 21.975)
MU9413/4/134 G_DS U9413/2/ix2093/B U9413/4/ix2099/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(18.69 21.715 18.82 21.975)
MU9413/4/135 G_DS U9413/4/ix2276/A U9413/4/136 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(19.87 21.715 20 22.015)
MU9413/4/136 U9413/2/ix2147/B U9413/4/136 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(20.45 21.715 20.58 22.015)
MU9413/4/137 U9413/4/ix2117/OUT wrData[13] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(21.63 21.715 21.76 21.975)
MU9413/4/138 G_DS U9413/2/ix2093/B U9413/4/ix2117/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(22.21 21.715 22.34 21.975)
MU9413/4/139 U9413/4/ix229/OUT U9413/3/ix2115/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(23.39 21.715 23.52 21.975)
MU9413/4/140 G_DS U9413/4/ix2117/OUT U9413/4/ix229/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(23.97 21.715 24.1 21.975)
MU9413/4/141 G_DS U9413/4/CLK U9413/4/144 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(25.15 21.715 25.28 22.015)
MU9413/4/142 U9413/4/145 U9413/4/144 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(25.73 21.715 25.86 22.015)
MU9413/4/143 U9413/4/146 U9413/3/ix217/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(26.82 21.715 26.95 22.105)
MU9413/4/144 U9413/4/148 U9413/4/145 U9413/4/146 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(27.335 21.715 27.465 22.105)
MU9413/4/145 U9413/4/149 U9413/4/148 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(28.425 21.715 28.555 22.015)
MU9413/4/146 U9413/4/150 U9413/4/144 U9413/4/148 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(29.515 21.715 29.645 22.105)
MU9413/4/147 G_DS U9413/4/CLB U9413/4/150 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(30.135 21.715 30.265 22.105)
MU9413/4/148 U9413/4/150 U9413/4/149 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(30.755 21.715 30.885 22.105)
MU9413/4/149 U9413/4/151 U9413/4/149 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(31.845 21.715 31.975 22.105)
MU9413/4/150 U9413/4/152 U9413/4/144 U9413/4/151 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(32.155 21.715 32.285 22.105)
MU9413/4/151 U9413/4/153 U9413/4/152 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(33.865 21.715 33.995 22.015)
MU9413/4/152 U9413/4/154 U9413/4/145 U9413/4/152 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(34.955 21.715 35.085 22.105)
MU9413/4/153 G_DS U9413/4/CLB U9413/4/154 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(35.535 21.715 35.665 22.105)
MU9413/4/154 U9413/4/154 U9413/4/153 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(36.115 21.715 36.245 22.015)
MU9413/4/155 wrData[13] U9413/4/154 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(37.205 21.715 37.335 22.015)
MU9413/4/156 U9413/4/reg_r_shiftReg_14_/QB U9413/4/153 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(38.295 21.715 38.425 22.015)
MU9413/4/157 G_DS U9413/4/CLK U9413/4/157 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(39.475 21.715 39.605 22.015)
MU9413/4/158 U9413/4/158 U9413/4/157 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(40.055 21.715 40.185 22.015)
MU9413/4/159 U9413/4/159 U9413/3/ix193/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(41.145 21.715 41.275 22.105)
MU9413/4/160 U9413/4/161 U9413/4/158 U9413/4/159 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(41.66 21.715 41.79 22.105)
MU9413/4/161 U9413/4/162 U9413/4/161 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(42.75 21.715 42.88 22.015)
MU9413/4/162 U9413/4/163 U9413/4/157 U9413/4/161 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(43.84 21.715 43.97 22.105)
MU9413/4/163 G_DS U9413/4/CLB U9413/4/163 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(44.46 21.715 44.59 22.105)
MU9413/4/164 U9413/4/163 U9413/4/162 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(45.08 21.715 45.21 22.105)
MU9413/4/165 U9413/4/164 U9413/4/162 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(46.17 21.715 46.3 22.105)
MU9413/4/166 U9413/4/165 U9413/4/157 U9413/4/164 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(46.48 21.715 46.61 22.105)
MU9413/4/167 U9413/4/166 U9413/4/165 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(48.19 21.715 48.32 22.015)
MU9413/4/168 U9413/4/167 U9413/4/158 U9413/4/165 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(49.28 21.715 49.41 22.105)
MU9413/4/169 G_DS U9413/4/CLB U9413/4/167 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(49.86 21.715 49.99 22.105)
MU9413/4/170 U9413/4/167 U9413/4/166 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(50.44 21.715 50.57 22.015)
MU9413/4/171 wrData[11] U9413/4/167 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(51.53 21.715 51.66 22.015)
MU9413/4/172 U9413/4/reg_r_shiftReg_12_/QB U9413/4/166 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(52.62 21.715 52.75 22.015)
MU9413/4/173 U9413/4/ix205/B wrData[11] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(53.8 21.715 53.93 21.975)
MU9413/4/174 G_DS U9413/2/ix2093/B U9413/4/ix205/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(54.38 21.715 54.51 21.975)
MU9413/4/175 U9413/4/ix205/OUT U9413/2/ix2127/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(55.56 21.715 55.69 21.975)
MU9413/4/176 G_DS U9413/4/ix205/B U9413/4/ix205/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(56.14 21.715 56.27 21.975)
MU9413/4/177 U9413/4/ix157/B wrData[7] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(57.32 21.715 57.45 21.975)
MU9413/4/178 G_DS U9413/2/ix2147/B U9413/4/ix157/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(57.9 21.715 58.03 21.975)
MU9413/4/179 U9413/reg_r_shiftReg_13_\Cross U9413/3/ix2151/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(59.08 21.715 59.21 21.975)
MU9413/4/180 G_DS U9413/4/ix157/B U9413/reg_r_shiftReg_13_\Cross G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(59.66 21.715 59.79 21.975)
MU9413/4/181 U9413/4/ix145/B wrData[6] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(60.84 21.715 60.97 21.975)
MU9413/4/182 G_DS U9413/2/ix2147/B U9413/4/ix145/B G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(61.42 21.715 61.55 21.975)
MU9413/4/183 U9413/4/ix145/OUT U9413/3/ix2157/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(62.6 21.715 62.73 21.975)
MU9413/4/184 G_DS U9413/4/ix145/B U9413/4/ix145/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(63.18 21.715 63.31 21.975)
MU9413/4/185 G_DS U9413/4/CLK U9413/4/188 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(64.36 21.715 64.49 22.015)
MU9413/4/186 U9413/4/189 U9413/4/188 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(64.94 21.715 65.07 22.015)
MU9413/4/187 U9413/4/190 U9413/3/ix133/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(66.03 21.715 66.16 22.105)
MU9413/4/188 U9413/4/192 U9413/4/189 U9413/4/190 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(66.545 21.715 66.675 22.105)
MU9413/4/189 U9413/4/193 U9413/4/192 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(67.635 21.715 67.765 22.015)
MU9413/4/190 U9413/4/194 U9413/4/188 U9413/4/192 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(68.725 21.715 68.855 22.105)
MU9413/4/191 G_DS U9413/4/CLB U9413/4/194 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(69.345 21.715 69.475 22.105)
MU9413/4/192 U9413/4/194 U9413/4/193 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(69.965 21.715 70.095 22.105)
MU9413/4/193 U9413/4/195 U9413/4/193 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(71.055 21.715 71.185 22.105)
MU9413/4/194 U9413/4/196 U9413/4/188 U9413/4/195 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(71.365 21.715 71.495 22.105)
MU9413/4/195 U9413/4/197 U9413/4/196 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(73.075 21.715 73.205 22.015)
MU9413/4/196 U9413/4/198 U9413/4/189 U9413/4/196 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(74.165 21.715 74.295 22.105)
MU9413/4/197 G_DS U9413/4/CLB U9413/4/198 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(74.745 21.715 74.875 22.105)
MU9413/4/198 U9413/4/198 U9413/4/197 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(75.325 21.715 75.455 22.015)
MU9413/4/199 wrData[6] U9413/4/198 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(76.415 21.715 76.545 22.015)
MU9413/4/200 U9413/4/reg_r_shiftReg_7_/QB U9413/4/197 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(77.505 21.715 77.635 22.015)
MU9413/4/201 G_DS U9413/4/CLK U9413/4/201 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(78.685 21.715 78.815 22.015)
MU9413/4/202 U9413/4/202 U9413/4/201 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(79.265 21.715 79.395 22.015)
MU9413/4/203 U9413/4/203 U9413/4/ix97/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(80.355 21.715 80.485 22.105)
MU9413/4/204 U9413/4/205 U9413/4/202 U9413/4/203 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(80.87 21.715 81 22.105)
MU9413/4/205 U9413/4/206 U9413/4/205 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(81.96 21.715 82.09 22.015)
MU9413/4/206 U9413/4/207 U9413/4/201 U9413/4/205 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(83.05 21.715 83.18 22.105)
MU9413/4/207 G_DS U9413/4/CLB U9413/4/207 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(83.67 21.715 83.8 22.105)
MU9413/4/208 U9413/4/207 U9413/4/206 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(84.29 21.715 84.42 22.105)
MU9413/4/209 U9413/4/208 U9413/4/206 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(85.38 21.715 85.51 22.105)
MU9413/4/210 U9413/4/209 U9413/4/201 U9413/4/208 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(85.69 21.715 85.82 22.105)
MU9413/4/211 U9413/4/210 U9413/4/209 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(87.4 21.715 87.53 22.015)
MU9413/4/212 U9413/4/211 U9413/4/202 U9413/4/209 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(88.49 21.715 88.62 22.105)
MU9413/4/213 G_DS U9413/4/CLB U9413/4/211 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(89.07 21.715 89.2 22.105)
MU9413/4/214 U9413/4/211 U9413/4/210 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(89.65 21.715 89.78 22.015)
MU9413/4/215 wrData[3] U9413/4/211 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(90.74 21.715 90.87 22.015)
MU9413/4/216 U9413/4/reg_r_shiftReg_4_/QB U9413/4/210 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(91.83 21.715 91.96 22.015)
MU9413/4/217 U9413/4/ix97/OUT U9413/3/ix2181/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(93.01 21.715 93.14 21.975)
MU9413/4/218 G_DS U9413/4/ix2183/OUT U9413/4/ix97/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(93.59 21.715 93.72 21.975)
MU9413/4/219 U9413/4/ix2183/OUT wrData[2] G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(94.77 21.715 94.9 21.975)
MU9413/4/220 G_DS U9413/2/ix2147/B U9413/4/ix2183/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(95.35 21.715 95.48 21.975)
MU9413/4/221 G_DS U9413/4/CLK U9413/4/220 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(96.53 21.715 96.66 22.015)
MU9413/4/222 U9413/4/221 U9413/4/220 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(97.11 21.715 97.24 22.015)
MU9413/4/223 U9413/4/222 U9413/4/ix1786/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(98.2 21.715 98.33 22.105)
MU9413/4/224 U9413/4/224 U9413/4/221 U9413/4/222 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(98.715 21.715 98.845 22.105)
MU9413/4/225 U9413/4/225 U9413/4/224 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(99.805 21.715 99.935 22.015)
MU9413/4/226 U9413/4/226 U9413/4/220 U9413/4/224 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(100.895 21.715 101.025 22.105)
MU9413/4/227 G_DS U9413/4/CLB U9413/4/226 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(101.515 21.715 101.645 22.105)
MU9413/4/228 U9413/4/226 U9413/4/225 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(102.135 21.715 102.265 22.105)
MU9413/4/229 U9413/4/227 U9413/4/225 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(103.225 21.715 103.355 22.105)
MU9413/4/230 U9413/4/228 U9413/4/220 U9413/4/227 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(103.535 21.715 103.665 22.105)
MU9413/4/231 U9413/4/229 U9413/4/228 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(105.245 21.715 105.375 22.015)
MU9413/4/232 U9413/4/230 U9413/4/221 U9413/4/228 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(106.335 21.715 106.465 22.105)
MU9413/4/233 G_DS U9413/4/CLB U9413/4/230 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(106.915 21.715 107.045 22.105)
MU9413/4/234 U9413/4/230 U9413/4/229 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(107.495 21.715 107.625 22.015)
MU9413/4/235 addr[8] U9413/4/230 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(108.585 21.715 108.715 22.015)
MU9413/4/236 U9413/4/reg_r_shiftReg_41_/QB U9413/4/229 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(109.675 21.715 109.805 22.015)
MU9413/4/237 G_DS U9413/SEL U9413/4/234 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(110.855 21.5 110.985 21.8)
MU9413/4/238 U9413/4/235 U9413/4/234 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(111.435 21.5 111.565 22.02)
MU9413/4/239 U9413/4/236 addr[7] U9413/4/235 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(112.015 21.5 112.145 22.02)
MU9413/4/240 U9413/4/238 addr[8] U9413/4/236 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(112.595 21.5 112.725 22.02)
MU9413/4/241 G_DS U9413/SEL U9413/4/238 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(113.175 21.5 113.305 22.02)
MU9413/4/242 U9413/4/ix1786/OUT U9413/4/236 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(113.755 21.715 113.885 22.015)
MU9413/4/243 G_DS U9413/SEL U9413/4/241 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(114.935 21.5 115.065 21.8)
MU9413/4/244 U9413/4/242 U9413/4/241 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(115.515 21.5 115.645 22.02)
MU9413/4/245 U9413/4/243 addr[8] U9413/4/242 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(116.095 21.5 116.225 22.02)
MU9413/4/246 U9413/4/244 addr[9] U9413/4/243 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(116.675 21.5 116.805 22.02)
MU9413/4/247 G_DS U9413/SEL U9413/4/244 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(117.255 21.5 117.385 22.02)
MU9413/4/248 U9413/4/DATA U9413/4/243 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(117.835 21.715 117.965 22.015)
MU9413/4/249 G_DS U9413/4/CLK U9413/4/245 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(119.015 21.715 119.145 22.015)
MU9413/4/250 U9413/4/246 U9413/4/245 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(119.595 21.715 119.725 22.015)
MU9413/4/251 U9413/4/247 U9413/4/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(120.685 21.715 120.815 22.105)
MU9413/4/252 U9413/4/248 U9413/4/246 U9413/4/247 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(121.2 21.715 121.33 22.105)
MU9413/4/253 U9413/4/249 U9413/4/248 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(122.29 21.715 122.42 22.015)
MU9413/4/254 U9413/4/250 U9413/4/245 U9413/4/248 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(123.38 21.715 123.51 22.105)
MU9413/4/255 G_DS U9413/4/CLB U9413/4/250 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(124 21.715 124.13 22.105)
MU9413/4/256 U9413/4/250 U9413/4/249 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(124.62 21.715 124.75 22.105)
MU9413/4/257 U9413/4/251 U9413/4/249 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(125.71 21.715 125.84 22.105)
MU9413/4/258 U9413/4/252 U9413/4/245 U9413/4/251 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(126.02 21.715 126.15 22.105)
MU9413/4/259 U9413/4/253 U9413/4/252 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(127.73 21.715 127.86 22.015)
MU9413/4/260 U9413/4/254 U9413/4/246 U9413/4/252 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(128.82 21.715 128.95 22.105)
MU9413/4/261 G_DS U9413/4/CLB U9413/4/254 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(129.4 21.715 129.53 22.105)
MU9413/4/262 U9413/4/254 U9413/4/253 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(129.98 21.715 130.11 22.015)
MU9413/4/263 addr[9] U9413/4/254 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(131.07 21.715 131.2 22.015)
MU9413/4/264 U9413/4/reg_r_shiftReg_42_/QB U9413/4/253 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(132.16 21.715 132.29 22.015)
MU9413/4/265 G_DS RST U9413/4/256 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(133.34 21.715 133.47 22.015)
MU9413/4/266 U9413/4/CLB U9413/4/256 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(133.92 21.715 134.05 22.015)
MU9413/4/267 G_DS RST U9413/4/257 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(135.1 21.715 135.23 22.015)
MU9413/4/268 U9413/4/CLB U9413/4/257 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(135.68 21.715 135.81 22.015)
MU9413/4/right_31/1 G_DG RST U9413/4/256 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(133.34 19.985 133.47 20.135)
MU9413/4/right_31/2 U9413/4/CLB U9413/4/256 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(133.92 19.985 134.05 20.135)
MU9413/4/right_30/1 G_DG RST U9413/4/257 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(135.1 19.985 135.23 20.135)
MU9413/4/right_30/2 U9413/4/CLB U9413/4/257 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(135.68 19.985 135.81 20.135)
MU9413/4/left_31/1 G_DG CLK U9413/4/2 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-98.32 19.985 -98.19 20.135)
MU9413/4/left_31/2 U9413/4/CLK U9413/4/2 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-97.74 19.985 -97.61 20.135)
MU9413/4/left_30/1 G_DG CLK U9413/4/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-96.56 19.985 -96.43 20.135)
MU9413/4/left_30/2 U9413/4/CLK U9413/4/3 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-95.98 19.985 -95.85 20.135)
MU9413/4/reg_r_shiftReg_42_/1 G_DG U9413/4/CLK U9413/4/245 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(119.015 19.985 119.145 20.135)
MU9413/4/reg_r_shiftReg_42_/2 U9413/4/246 U9413/4/245 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(119.595 19.985 119.725 20.135)
MU9413/4/reg_r_shiftReg_42_/3 U9413/4/reg_r_shiftReg_42_/4 U9413/4/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(120.685 19.985 120.815 20.135)
MU9413/4/reg_r_shiftReg_42_/4 U9413/4/248 U9413/4/245 U9413/4/reg_r_shiftReg_42_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(121.2 19.985 121.33 20.135)
MU9413/4/reg_r_shiftReg_42_/5 U9413/4/249 U9413/4/248 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(122.29 19.985 122.42 20.135)
MU9413/4/reg_r_shiftReg_42_/6 U9413/4/reg_r_shiftReg_42_/7 U9413/4/CLB U9413/4/248 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(123.66 19.985 123.79 20.135)
MU9413/4/reg_r_shiftReg_42_/7 U9413/4/reg_r_shiftReg_42_/8 U9413/4/249 U9413/4/reg_r_shiftReg_42_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(124.14 19.985 124.27 20.135)
MU9413/4/reg_r_shiftReg_42_/8 G_DG U9413/4/246 U9413/4/reg_r_shiftReg_42_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(124.62 19.985 124.75 20.135)
MU9413/4/reg_r_shiftReg_42_/9 U9413/4/reg_r_shiftReg_42_/9 U9413/4/249 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(125.71 19.985 125.84 20.135)
MU9413/4/reg_r_shiftReg_42_/10 U9413/4/reg_r_shiftReg_42_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_42_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(126.22 19.985 126.35 20.135)
MU9413/4/reg_r_shiftReg_42_/11 U9413/4/252 U9413/4/246 U9413/4/reg_r_shiftReg_42_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(126.64 19.985 126.77 20.135)
MU9413/4/reg_r_shiftReg_42_/12 U9413/4/253 U9413/4/252 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(127.73 19.985 127.86 20.135)
MU9413/4/reg_r_shiftReg_42_/13 U9413/4/254 U9413/4/245 U9413/4/252 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(129.09 19.985 129.22 20.135)
MU9413/4/reg_r_shiftReg_42_/14 U9413/4/reg_r_shiftReg_42_/14 U9413/4/CLB U9413/4/254 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(129.67 19.985 129.8 20.135)
MU9413/4/reg_r_shiftReg_42_/15 G_DG U9413/4/253 U9413/4/reg_r_shiftReg_42_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(129.98 19.985 130.11 20.135)
MU9413/4/reg_r_shiftReg_42_/16 addr[9] U9413/4/254 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(131.07 19.985 131.2 20.135)
MU9413/4/reg_r_shiftReg_42_/17 U9413/4/reg_r_shiftReg_42_/QB U9413/4/253 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(132.16 19.985 132.29 20.135)
MU9413/4/ix1796/1 G_DG U9413/SEL U9413/4/241 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(114.935 19.985 115.065 20.135)
MU9413/4/ix1796/2 U9413/4/ix1796/3 U9413/4/241 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(115.515 19.985 115.645 20.135)
MU9413/4/ix1796/3 U9413/4/243 addr[9] U9413/4/ix1796/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(116.095 19.985 116.225 20.135)
MU9413/4/ix1796/4 U9413/4/ix1796/5 addr[8] U9413/4/243 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(116.675 19.985 116.805 20.135)
MU9413/4/ix1796/5 G_DG U9413/SEL U9413/4/ix1796/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(117.255 19.985 117.385 20.135)
MU9413/4/ix1796/6 U9413/4/DATA U9413/4/243 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(117.835 19.985 117.965 20.135)
MU9413/4/ix1786/1 G_DG U9413/SEL U9413/4/234 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(110.855 19.985 110.985 20.135)
MU9413/4/ix1786/2 U9413/4/ix1786/3 U9413/4/234 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(111.435 19.985 111.565 20.135)
MU9413/4/ix1786/3 U9413/4/236 addr[8] U9413/4/ix1786/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(112.015 19.985 112.145 20.135)
MU9413/4/ix1786/4 U9413/4/ix1786/5 addr[7] U9413/4/236 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(112.595 19.985 112.725 20.135)
MU9413/4/ix1786/5 G_DG U9413/SEL U9413/4/ix1786/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(113.175 19.985 113.305 20.135)
MU9413/4/ix1786/6 U9413/4/ix1786/OUT U9413/4/236 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(113.755 19.985 113.885 20.135)
MU9413/4/reg_r_shiftReg_41_/1 G_DG U9413/4/CLK U9413/4/220 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(96.53 19.985 96.66 20.135)
MU9413/4/reg_r_shiftReg_41_/2 U9413/4/221 U9413/4/220 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(97.11 19.985 97.24 20.135)
MU9413/4/reg_r_shiftReg_41_/3 U9413/4/reg_r_shiftReg_41_/4 U9413/4/ix1786/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(98.2 19.985 98.33 20.135)
MU9413/4/reg_r_shiftReg_41_/4 U9413/4/224 U9413/4/220 U9413/4/reg_r_shiftReg_41_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(98.715 19.985 98.845 20.135)
MU9413/4/reg_r_shiftReg_41_/5 U9413/4/225 U9413/4/224 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(99.805 19.985 99.935 20.135)
MU9413/4/reg_r_shiftReg_41_/6 U9413/4/reg_r_shiftReg_41_/7 U9413/4/CLB U9413/4/224 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(101.175 19.985 101.305 20.135)
MU9413/4/reg_r_shiftReg_41_/7 U9413/4/reg_r_shiftReg_41_/8 U9413/4/225 U9413/4/reg_r_shiftReg_41_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(101.655 19.985 101.785 20.135)
MU9413/4/reg_r_shiftReg_41_/8 G_DG U9413/4/221 U9413/4/reg_r_shiftReg_41_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(102.135 19.985 102.265 20.135)
MU9413/4/reg_r_shiftReg_41_/9 U9413/4/reg_r_shiftReg_41_/9 U9413/4/225 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(103.225 19.985 103.355 20.135)
MU9413/4/reg_r_shiftReg_41_/10 U9413/4/reg_r_shiftReg_41_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_41_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(103.735 19.985 103.865 20.135)
MU9413/4/reg_r_shiftReg_41_/11 U9413/4/228 U9413/4/221 U9413/4/reg_r_shiftReg_41_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(104.155 19.985 104.285 20.135)
MU9413/4/reg_r_shiftReg_41_/12 U9413/4/229 U9413/4/228 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(105.245 19.985 105.375 20.135)
MU9413/4/reg_r_shiftReg_41_/13 U9413/4/230 U9413/4/220 U9413/4/228 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(106.605 19.985 106.735 20.135)
MU9413/4/reg_r_shiftReg_41_/14 U9413/4/reg_r_shiftReg_41_/14 U9413/4/CLB U9413/4/230 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(107.185 19.985 107.315 20.135)
MU9413/4/reg_r_shiftReg_41_/15 G_DG U9413/4/229 U9413/4/reg_r_shiftReg_41_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(107.495 19.985 107.625 20.135)
MU9413/4/reg_r_shiftReg_41_/16 addr[8] U9413/4/230 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(108.585 19.985 108.715 20.135)
MU9413/4/reg_r_shiftReg_41_/17 U9413/4/reg_r_shiftReg_41_/QB U9413/4/229 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(109.675 19.985 109.805 20.135)
MU9413/4/ix2183/1 U9413/4/ix2183/1 wrData[2] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(94.77 19.985 94.9 20.135)
MU9413/4/ix2183/2 U9413/4/ix2183/OUT U9413/2/ix2147/B U9413/4/ix2183/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(95.35 19.985 95.48 20.135)
MU9413/4/ix97/1 U9413/4/ix97/1 U9413/3/ix2181/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(93.01 19.985 93.14 20.135)
MU9413/4/ix97/2 U9413/4/ix97/OUT U9413/4/ix2183/OUT U9413/4/ix97/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(93.59 19.985 93.72 20.135)
MU9413/4/reg_r_shiftReg_4_/1 G_DG U9413/4/CLK U9413/4/201 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(78.685 19.985 78.815 20.135)
MU9413/4/reg_r_shiftReg_4_/2 U9413/4/202 U9413/4/201 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(79.265 19.985 79.395 20.135)
MU9413/4/reg_r_shiftReg_4_/3 U9413/4/reg_r_shiftReg_4_/4 U9413/4/ix97/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(80.355 19.985 80.485 20.135)
MU9413/4/reg_r_shiftReg_4_/4 U9413/4/205 U9413/4/201 U9413/4/reg_r_shiftReg_4_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(80.87 19.985 81 20.135)
MU9413/4/reg_r_shiftReg_4_/5 U9413/4/206 U9413/4/205 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(81.96 19.985 82.09 20.135)
MU9413/4/reg_r_shiftReg_4_/6 U9413/4/reg_r_shiftReg_4_/7 U9413/4/CLB U9413/4/205 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(83.33 19.985 83.46 20.135)
MU9413/4/reg_r_shiftReg_4_/7 U9413/4/reg_r_shiftReg_4_/8 U9413/4/206 U9413/4/reg_r_shiftReg_4_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(83.81 19.985 83.94 20.135)
MU9413/4/reg_r_shiftReg_4_/8 G_DG U9413/4/202 U9413/4/reg_r_shiftReg_4_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(84.29 19.985 84.42 20.135)
MU9413/4/reg_r_shiftReg_4_/9 U9413/4/reg_r_shiftReg_4_/9 U9413/4/206 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(85.38 19.985 85.51 20.135)
MU9413/4/reg_r_shiftReg_4_/10 U9413/4/reg_r_shiftReg_4_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_4_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(85.89 19.985 86.02 20.135)
MU9413/4/reg_r_shiftReg_4_/11 U9413/4/209 U9413/4/202 U9413/4/reg_r_shiftReg_4_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(86.31 19.985 86.44 20.135)
MU9413/4/reg_r_shiftReg_4_/12 U9413/4/210 U9413/4/209 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(87.4 19.985 87.53 20.135)
MU9413/4/reg_r_shiftReg_4_/13 U9413/4/211 U9413/4/201 U9413/4/209 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(88.76 19.985 88.89 20.135)
MU9413/4/reg_r_shiftReg_4_/14 U9413/4/reg_r_shiftReg_4_/14 U9413/4/CLB U9413/4/211 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(89.34 19.985 89.47 20.135)
MU9413/4/reg_r_shiftReg_4_/15 G_DG U9413/4/210 U9413/4/reg_r_shiftReg_4_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(89.65 19.985 89.78 20.135)
MU9413/4/reg_r_shiftReg_4_/16 wrData[3] U9413/4/211 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(90.74 19.985 90.87 20.135)
MU9413/4/reg_r_shiftReg_4_/17 U9413/4/reg_r_shiftReg_4_/QB U9413/4/210 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(91.83 19.985 91.96 20.135)
MU9413/4/reg_r_shiftReg_7_/1 G_DG U9413/4/CLK U9413/4/188 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(64.36 19.985 64.49 20.135)
MU9413/4/reg_r_shiftReg_7_/2 U9413/4/189 U9413/4/188 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(64.94 19.985 65.07 20.135)
MU9413/4/reg_r_shiftReg_7_/3 U9413/4/reg_r_shiftReg_7_/4 U9413/3/ix133/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(66.03 19.985 66.16 20.135)
MU9413/4/reg_r_shiftReg_7_/4 U9413/4/192 U9413/4/188 U9413/4/reg_r_shiftReg_7_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(66.545 19.985 66.675 20.135)
MU9413/4/reg_r_shiftReg_7_/5 U9413/4/193 U9413/4/192 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(67.635 19.985 67.765 20.135)
MU9413/4/reg_r_shiftReg_7_/6 U9413/4/reg_r_shiftReg_7_/7 U9413/4/CLB U9413/4/192 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(69.005 19.985 69.135 20.135)
MU9413/4/reg_r_shiftReg_7_/7 U9413/4/reg_r_shiftReg_7_/8 U9413/4/193 U9413/4/reg_r_shiftReg_7_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(69.485 19.985 69.615 20.135)
MU9413/4/reg_r_shiftReg_7_/8 G_DG U9413/4/189 U9413/4/reg_r_shiftReg_7_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(69.965 19.985 70.095 20.135)
MU9413/4/reg_r_shiftReg_7_/9 U9413/4/reg_r_shiftReg_7_/9 U9413/4/193 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(71.055 19.985 71.185 20.135)
MU9413/4/reg_r_shiftReg_7_/10 U9413/4/reg_r_shiftReg_7_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_7_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(71.565 19.985 71.695 20.135)
MU9413/4/reg_r_shiftReg_7_/11 U9413/4/196 U9413/4/189 U9413/4/reg_r_shiftReg_7_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(71.985 19.985 72.115 20.135)
MU9413/4/reg_r_shiftReg_7_/12 U9413/4/197 U9413/4/196 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(73.075 19.985 73.205 20.135)
MU9413/4/reg_r_shiftReg_7_/13 U9413/4/198 U9413/4/188 U9413/4/196 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(74.435 19.985 74.565 20.135)
MU9413/4/reg_r_shiftReg_7_/14 U9413/4/reg_r_shiftReg_7_/14 U9413/4/CLB U9413/4/198 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(75.015 19.985 75.145 20.135)
MU9413/4/reg_r_shiftReg_7_/15 G_DG U9413/4/197 U9413/4/reg_r_shiftReg_7_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(75.325 19.985 75.455 20.135)
MU9413/4/reg_r_shiftReg_7_/16 wrData[6] U9413/4/198 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(76.415 19.985 76.545 20.135)
MU9413/4/reg_r_shiftReg_7_/17 U9413/4/reg_r_shiftReg_7_/QB U9413/4/197 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(77.505 19.985 77.635 20.135)
MU9413/4/ix145/1 U9413/4/ix145/1 U9413/3/ix2157/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(62.6 19.985 62.73 20.135)
MU9413/4/ix145/2 U9413/4/ix145/OUT U9413/4/ix145/B U9413/4/ix145/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(63.18 19.985 63.31 20.135)
MU9413/4/ix2159/1 U9413/4/ix2159/1 wrData[6] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(60.84 19.985 60.97 20.135)
MU9413/4/ix2159/2 U9413/4/ix145/B U9413/2/ix2147/B U9413/4/ix2159/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(61.42 19.985 61.55 20.135)
MU9413/4/ix157/1 U9413/4/ix157/1 U9413/3/ix2151/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(59.08 19.985 59.21 20.135)
MU9413/4/ix157/2 U9413/reg_r_shiftReg_13_\Cross U9413/4/ix157/B U9413/4/ix157/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(59.66 19.985 59.79 20.135)
MU9413/4/ix2153/1 U9413/4/ix2153/1 wrData[7] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(57.32 19.985 57.45 20.135)
MU9413/4/ix2153/2 U9413/4/ix157/B U9413/2/ix2147/B U9413/4/ix2153/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(57.9 19.985 58.03 20.135)
MU9413/4/ix205/1 U9413/4/ix205/1 U9413/2/ix2127/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(55.56 19.985 55.69 20.135)
MU9413/4/ix205/2 U9413/4/ix205/OUT U9413/4/ix205/B U9413/4/ix205/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(56.14 19.985 56.27 20.135)
MU9413/4/ix2129/1 U9413/4/ix2129/1 wrData[11] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(53.8 19.985 53.93 20.135)
MU9413/4/ix2129/2 U9413/4/ix205/B U9413/2/ix2093/B U9413/4/ix2129/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(54.38 19.985 54.51 20.135)
MU9413/4/reg_r_shiftReg_12_/1 G_DG U9413/4/CLK U9413/4/157 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(39.475 19.985 39.605 20.135)
MU9413/4/reg_r_shiftReg_12_/2 U9413/4/158 U9413/4/157 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(40.055 19.985 40.185 20.135)
MU9413/4/reg_r_shiftReg_12_/3 U9413/4/reg_r_shiftReg_12_/4 U9413/3/ix193/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(41.145 19.985 41.275 20.135)
MU9413/4/reg_r_shiftReg_12_/4 U9413/4/161 U9413/4/157 U9413/4/reg_r_shiftReg_12_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(41.66 19.985 41.79 20.135)
MU9413/4/reg_r_shiftReg_12_/5 U9413/4/162 U9413/4/161 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(42.75 19.985 42.88 20.135)
MU9413/4/reg_r_shiftReg_12_/6 U9413/4/reg_r_shiftReg_12_/7 U9413/4/CLB U9413/4/161 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(44.12 19.985 44.25 20.135)
MU9413/4/reg_r_shiftReg_12_/7 U9413/4/reg_r_shiftReg_12_/8 U9413/4/162 U9413/4/reg_r_shiftReg_12_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(44.6 19.985 44.73 20.135)
MU9413/4/reg_r_shiftReg_12_/8 G_DG U9413/4/158 U9413/4/reg_r_shiftReg_12_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(45.08 19.985 45.21 20.135)
MU9413/4/reg_r_shiftReg_12_/9 U9413/4/reg_r_shiftReg_12_/9 U9413/4/162 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(46.17 19.985 46.3 20.135)
MU9413/4/reg_r_shiftReg_12_/10 U9413/4/reg_r_shiftReg_12_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_12_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(46.68 19.985 46.81 20.135)
MU9413/4/reg_r_shiftReg_12_/11 U9413/4/165 U9413/4/158 U9413/4/reg_r_shiftReg_12_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(47.1 19.985 47.23 20.135)
MU9413/4/reg_r_shiftReg_12_/12 U9413/4/166 U9413/4/165 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(48.19 19.985 48.32 20.135)
MU9413/4/reg_r_shiftReg_12_/13 U9413/4/167 U9413/4/157 U9413/4/165 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(49.55 19.985 49.68 20.135)
MU9413/4/reg_r_shiftReg_12_/14 U9413/4/reg_r_shiftReg_12_/14 U9413/4/CLB U9413/4/167 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(50.13 19.985 50.26 20.135)
MU9413/4/reg_r_shiftReg_12_/15 G_DG U9413/4/166 U9413/4/reg_r_shiftReg_12_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(50.44 19.985 50.57 20.135)
MU9413/4/reg_r_shiftReg_12_/16 wrData[11] U9413/4/167 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(51.53 19.985 51.66 20.135)
MU9413/4/reg_r_shiftReg_12_/17 U9413/4/reg_r_shiftReg_12_/QB U9413/4/166 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(52.62 19.985 52.75 20.135)
MU9413/4/reg_r_shiftReg_14_/1 G_DG U9413/4/CLK U9413/4/144 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(25.15 19.985 25.28 20.135)
MU9413/4/reg_r_shiftReg_14_/2 U9413/4/145 U9413/4/144 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(25.73 19.985 25.86 20.135)
MU9413/4/reg_r_shiftReg_14_/3 U9413/4/reg_r_shiftReg_14_/4 U9413/3/ix217/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(26.82 19.985 26.95 20.135)
MU9413/4/reg_r_shiftReg_14_/4 U9413/4/148 U9413/4/144 U9413/4/reg_r_shiftReg_14_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(27.335 19.985 27.465 20.135)
MU9413/4/reg_r_shiftReg_14_/5 U9413/4/149 U9413/4/148 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(28.425 19.985 28.555 20.135)
MU9413/4/reg_r_shiftReg_14_/6 U9413/4/reg_r_shiftReg_14_/7 U9413/4/CLB U9413/4/148 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(29.795 19.985 29.925 20.135)
MU9413/4/reg_r_shiftReg_14_/7 U9413/4/reg_r_shiftReg_14_/8 U9413/4/149 U9413/4/reg_r_shiftReg_14_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(30.275 19.985 30.405 20.135)
MU9413/4/reg_r_shiftReg_14_/8 G_DG U9413/4/145 U9413/4/reg_r_shiftReg_14_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(30.755 19.985 30.885 20.135)
MU9413/4/reg_r_shiftReg_14_/9 U9413/4/reg_r_shiftReg_14_/9 U9413/4/149 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(31.845 19.985 31.975 20.135)
MU9413/4/reg_r_shiftReg_14_/10 U9413/4/reg_r_shiftReg_14_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_14_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(32.355 19.985 32.485 20.135)
MU9413/4/reg_r_shiftReg_14_/11 U9413/4/152 U9413/4/145 U9413/4/reg_r_shiftReg_14_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(32.775 19.985 32.905 20.135)
MU9413/4/reg_r_shiftReg_14_/12 U9413/4/153 U9413/4/152 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(33.865 19.985 33.995 20.135)
MU9413/4/reg_r_shiftReg_14_/13 U9413/4/154 U9413/4/144 U9413/4/152 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(35.225 19.985 35.355 20.135)
MU9413/4/reg_r_shiftReg_14_/14 U9413/4/reg_r_shiftReg_14_/14 U9413/4/CLB U9413/4/154 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(35.805 19.985 35.935 20.135)
MU9413/4/reg_r_shiftReg_14_/15 G_DG U9413/4/153 U9413/4/reg_r_shiftReg_14_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(36.115 19.985 36.245 20.135)
MU9413/4/reg_r_shiftReg_14_/16 wrData[13] U9413/4/154 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(37.205 19.985 37.335 20.135)
MU9413/4/reg_r_shiftReg_14_/17 U9413/4/reg_r_shiftReg_14_/QB U9413/4/153 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(38.295 19.985 38.425 20.135)
MU9413/4/ix229/1 U9413/4/ix229/1 U9413/3/ix2115/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(23.39 19.985 23.52 20.135)
MU9413/4/ix229/2 U9413/4/ix229/OUT U9413/4/ix2117/OUT U9413/4/ix229/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(23.97 19.985 24.1 20.135)
MU9413/4/ix2117/1 U9413/4/ix2117/1 wrData[13] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(21.63 19.985 21.76 20.135)
MU9413/4/ix2117/2 U9413/4/ix2117/OUT U9413/2/ix2093/B U9413/4/ix2117/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(22.21 19.985 22.34 20.135)
MU9413/4/ix2276/1 G_DG U9413/4/ix2276/A U9413/4/136 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(19.87 19.985 20 20.135)
MU9413/4/ix2276/2 U9413/2/ix2147/B U9413/4/136 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(20.45 19.985 20.58 20.135)
MU9413/4/ix2099/1 U9413/4/ix2099/1 wrData[16] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(18.11 19.985 18.24 20.135)
MU9413/4/ix2099/2 U9413/4/ix2099/OUT U9413/2/ix2093/B U9413/4/ix2099/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(18.69 19.985 18.82 20.135)
MU9413/4/ix2278/1 G_DG U9413/4/ix2276/A U9413/4/130 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(16.35 19.985 16.48 20.135)
MU9413/4/ix2278/2 U9413/2/ix2093/B U9413/4/130 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(16.93 19.985 17.06 20.135)
MU9413/4/ix265/1 U9413/4/ix265/1 U9413/3/ix2097/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(14.59 19.985 14.72 20.135)
MU9413/4/ix265/2 U9413/4/ix265/OUT U9413/4/ix2099/OUT U9413/4/ix265/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(15.17 19.985 15.3 20.135)
MU9413/4/reg_r_shiftReg_18_/1 G_DG U9413/4/CLK U9413/4/113 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(0.265 19.985 0.395 20.135)
MU9413/4/reg_r_shiftReg_18_/2 U9413/4/114 U9413/4/113 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(0.845 19.985 0.975 20.135)
MU9413/4/reg_r_shiftReg_18_/3 U9413/4/reg_r_shiftReg_18_/4 U9413/4/ix265/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(1.935 19.985 2.065 20.135)
MU9413/4/reg_r_shiftReg_18_/4 U9413/4/117 U9413/4/113 U9413/4/reg_r_shiftReg_18_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(2.45 19.985 2.58 20.135)
MU9413/4/reg_r_shiftReg_18_/5 U9413/4/118 U9413/4/117 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(3.54 19.985 3.67 20.135)
MU9413/4/reg_r_shiftReg_18_/6 U9413/4/reg_r_shiftReg_18_/7 U9413/4/CLB U9413/4/117 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(4.91 19.985 5.04 20.135)
MU9413/4/reg_r_shiftReg_18_/7 U9413/4/reg_r_shiftReg_18_/8 U9413/4/118 U9413/4/reg_r_shiftReg_18_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(5.39 19.985 5.52 20.135)
MU9413/4/reg_r_shiftReg_18_/8 G_DG U9413/4/114 U9413/4/reg_r_shiftReg_18_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(5.87 19.985 6 20.135)
MU9413/4/reg_r_shiftReg_18_/9 U9413/4/reg_r_shiftReg_18_/9 U9413/4/118 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(6.96 19.985 7.09 20.135)
MU9413/4/reg_r_shiftReg_18_/10 U9413/4/reg_r_shiftReg_18_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_18_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(7.47 19.985 7.6 20.135)
MU9413/4/reg_r_shiftReg_18_/11 U9413/4/121 U9413/4/114 U9413/4/reg_r_shiftReg_18_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(7.89 19.985 8.02 20.135)
MU9413/4/reg_r_shiftReg_18_/12 U9413/4/122 U9413/4/121 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(8.98 19.985 9.11 20.135)
MU9413/4/reg_r_shiftReg_18_/13 U9413/4/123 U9413/4/113 U9413/4/121 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(10.34 19.985 10.47 20.135)
MU9413/4/reg_r_shiftReg_18_/14 U9413/4/reg_r_shiftReg_18_/14 U9413/4/CLB U9413/4/123 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(10.92 19.985 11.05 20.135)
MU9413/4/reg_r_shiftReg_18_/15 G_DG U9413/4/122 U9413/4/reg_r_shiftReg_18_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(11.23 19.985 11.36 20.135)
MU9413/4/reg_r_shiftReg_18_/16 wrData[17] U9413/4/123 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(12.32 19.985 12.45 20.135)
MU9413/4/reg_r_shiftReg_18_/17 U9413/4/reg_r_shiftReg_18_/QB U9413/4/122 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(13.41 19.985 13.54 20.135)
MU9413/4/ix2251/1 U9413/4/ix2251/1 U9413/4/ix2251/A G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-1.495 19.985 -1.365 20.135)
MU9413/4/ix2251/2 U9413/reg_r_shiftReg_21_\Cross U9413/2/ix2021/B U9413/4/ix2251/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-0.915 19.985 -0.785 20.135)
MU9413/4/ix2280/1 G_DG U9413/4/ix2276/A U9413/4/108 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-3.255 19.985 -3.125 20.135)
MU9413/4/ix2280/2 U9413/2/ix2045/B U9413/4/108 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-2.675 19.985 -2.545 20.135)
MU9413/4/ix2282/1 G_DG U9413/4/ix2276/A U9413/4/105 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-5.015 19.985 -4.885 20.135)
MU9413/4/ix2282/2 U9413/2/ix2021/B U9413/4/105 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-4.435 19.985 -4.305 20.135)
MU9413/4/ix2288/1 U9413/2/ix2121/D ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-6.775 19.985 -6.645 20.135)
MU9413/4/ix2288/2 G_DG U9413/4/ix2270/OUT U9413/2/ix2121/D G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-6.195 19.985 -6.065 20.135)
MU9413/4/ix2286/1 U9413/2/ix2067/D ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-8.535 19.985 -8.405 20.135)
MU9413/4/ix2286/2 G_DG U9413/4/ix2270/OUT U9413/2/ix2067/D G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-7.955 19.985 -7.825 20.135)
MU9413/4/ix2075/1 U9413/4/ix2075/1 wrData[20] G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-10.295 19.985 -10.165 20.135)
MU9413/4/ix2075/2 U9413/4/ix2075/OUT U9413/2/ix2045/B U9413/4/ix2075/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-9.715 19.985 -9.585 20.135)
MU9413/4/ix313/1 U9413/4/ix313/1 U9413/3/ix2073/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-12.055 19.985 -11.925 20.135)
MU9413/4/ix313/2 U9413/4/ix313/OUT U9413/4/ix2075/OUT U9413/4/ix313/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-11.475 19.985 -11.345 20.135)
MU9413/4/ix2290/1 G_DG U9413/3/ix2292/A U9413/4/88 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-13.815 19.985 -13.685 20.135)
MU9413/4/ix2290/2 U9413/2/ix2019/B U9413/4/88 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-13.235 19.985 -13.105 20.135)
MU9413/4/reg_r_shiftReg_22_/1 G_DG U9413/4/CLK U9413/4/74 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-28.14 19.985 -28.01 20.135)
MU9413/4/reg_r_shiftReg_22_/2 U9413/4/75 U9413/4/74 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-27.56 19.985 -27.43 20.135)
MU9413/4/reg_r_shiftReg_22_/3 U9413/4/reg_r_shiftReg_22_/4 U9413/4/ix313/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-26.47 19.985 -26.34 20.135)
MU9413/4/reg_r_shiftReg_22_/4 U9413/4/78 U9413/4/74 U9413/4/reg_r_shiftReg_22_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-25.955 19.985 -25.825 20.135)
MU9413/4/reg_r_shiftReg_22_/5 U9413/4/79 U9413/4/78 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-24.865 19.985 -24.735 20.135)
MU9413/4/reg_r_shiftReg_22_/6 U9413/4/reg_r_shiftReg_22_/7 U9413/4/CLB U9413/4/78 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-23.495 19.985 -23.365 20.135)
MU9413/4/reg_r_shiftReg_22_/7 U9413/4/reg_r_shiftReg_22_/8 U9413/4/79 U9413/4/reg_r_shiftReg_22_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-23.015 19.985 -22.885 20.135)
MU9413/4/reg_r_shiftReg_22_/8 G_DG U9413/4/75 U9413/4/reg_r_shiftReg_22_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-22.535 19.985 -22.405 20.135)
MU9413/4/reg_r_shiftReg_22_/9 U9413/4/reg_r_shiftReg_22_/9 U9413/4/79 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-21.445 19.985 -21.315 20.135)
MU9413/4/reg_r_shiftReg_22_/10 U9413/4/reg_r_shiftReg_22_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_22_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-20.935 19.985 -20.805 20.135)
MU9413/4/reg_r_shiftReg_22_/11 U9413/4/82 U9413/4/75 U9413/4/reg_r_shiftReg_22_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-20.515 19.985 -20.385 20.135)
MU9413/4/reg_r_shiftReg_22_/12 U9413/4/83 U9413/4/82 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-19.425 19.985 -19.295 20.135)
MU9413/4/reg_r_shiftReg_22_/13 U9413/4/84 U9413/4/74 U9413/4/82 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-18.065 19.985 -17.935 20.135)
MU9413/4/reg_r_shiftReg_22_/14 U9413/4/reg_r_shiftReg_22_/14 U9413/4/CLB U9413/4/84 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-17.485 19.985 -17.355 20.135)
MU9413/4/reg_r_shiftReg_22_/15 G_DG U9413/4/83 U9413/4/reg_r_shiftReg_22_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-17.175 19.985 -17.045 20.135)
MU9413/4/reg_r_shiftReg_22_/16 wrData[21] U9413/4/84 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-16.085 19.985 -15.955 20.135)
MU9413/4/reg_r_shiftReg_22_/17 U9413/4/reg_r_shiftReg_22_/QB U9413/4/83 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-14.995 19.985 -14.865 20.135)
MU9413/4/ix2270/1 G_DG U9413/4/ix2270/A U9413/4/72 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-29.9 19.985 -29.77 20.135)
MU9413/4/ix2270/2 U9413/4/ix2270/OUT U9413/4/72 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-29.32 19.985 -29.19 20.135)
MU9413/4/ix2284/1 U9413/2/ix2019/D ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-31.66 19.985 -31.53 20.135)
MU9413/4/ix2284/2 G_DG U9413/4/ix2270/OUT U9413/2/ix2019/D G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-31.08 19.985 -30.95 20.135)
MU9413/4/reg_r_shiftReg_25_/1 G_DG U9413/4/CLK U9413/4/54 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-45.985 19.985 -45.855 20.135)
MU9413/4/reg_r_shiftReg_25_/2 U9413/4/55 U9413/4/54 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-45.405 19.985 -45.275 20.135)
MU9413/4/reg_r_shiftReg_25_/3 U9413/4/reg_r_shiftReg_25_/4 U9413/3/ix349/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-44.315 19.985 -44.185 20.135)
MU9413/4/reg_r_shiftReg_25_/4 U9413/4/58 U9413/4/54 U9413/4/reg_r_shiftReg_25_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-43.8 19.985 -43.67 20.135)
MU9413/4/reg_r_shiftReg_25_/5 U9413/4/59 U9413/4/58 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-42.71 19.985 -42.58 20.135)
MU9413/4/reg_r_shiftReg_25_/6 U9413/4/reg_r_shiftReg_25_/7 U9413/4/CLB U9413/4/58 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-41.34 19.985 -41.21 20.135)
MU9413/4/reg_r_shiftReg_25_/7 U9413/4/reg_r_shiftReg_25_/8 U9413/4/59 U9413/4/reg_r_shiftReg_25_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-40.86 19.985 -40.73 20.135)
MU9413/4/reg_r_shiftReg_25_/8 G_DG U9413/4/55 U9413/4/reg_r_shiftReg_25_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-40.38 19.985 -40.25 20.135)
MU9413/4/reg_r_shiftReg_25_/9 U9413/4/reg_r_shiftReg_25_/9 U9413/4/59 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-39.29 19.985 -39.16 20.135)
MU9413/4/reg_r_shiftReg_25_/10 U9413/4/reg_r_shiftReg_25_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_25_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-38.78 19.985 -38.65 20.135)
MU9413/4/reg_r_shiftReg_25_/11 U9413/4/62 U9413/4/55 U9413/4/reg_r_shiftReg_25_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-38.36 19.985 -38.23 20.135)
MU9413/4/reg_r_shiftReg_25_/12 U9413/4/63 U9413/4/62 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-37.27 19.985 -37.14 20.135)
MU9413/4/reg_r_shiftReg_25_/13 U9413/4/64 U9413/4/54 U9413/4/62 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-35.91 19.985 -35.78 20.135)
MU9413/4/reg_r_shiftReg_25_/14 U9413/4/reg_r_shiftReg_25_/14 U9413/4/CLB U9413/4/64 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-35.33 19.985 -35.2 20.135)
MU9413/4/reg_r_shiftReg_25_/15 G_DG U9413/4/63 U9413/4/reg_r_shiftReg_25_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-35.02 19.985 -34.89 20.135)
MU9413/4/reg_r_shiftReg_25_/16 wrData[24] U9413/4/64 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-33.93 19.985 -33.8 20.135)
MU9413/4/reg_r_shiftReg_25_/17 U9413/4/reg_r_shiftReg_25_/QB U9413/4/63 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-32.84 19.985 -32.71 20.135)
MU9413/4/reg_r_shiftReg_28_/1 G_DG U9413/4/CLK U9413/4/41 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-60.31 19.985 -60.18 20.135)
MU9413/4/reg_r_shiftReg_28_/2 U9413/4/42 U9413/4/41 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-59.73 19.985 -59.6 20.135)
MU9413/4/reg_r_shiftReg_28_/3 U9413/4/reg_r_shiftReg_28_/4 U9413/3/ix385/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-58.64 19.985 -58.51 20.135)
MU9413/4/reg_r_shiftReg_28_/4 U9413/4/45 U9413/4/41 U9413/4/reg_r_shiftReg_28_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-58.125 19.985 -57.995 20.135)
MU9413/4/reg_r_shiftReg_28_/5 U9413/4/46 U9413/4/45 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-57.035 19.985 -56.905 20.135)
MU9413/4/reg_r_shiftReg_28_/6 U9413/4/reg_r_shiftReg_28_/7 U9413/4/CLB U9413/4/45 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-55.665 19.985 -55.535 20.135)
MU9413/4/reg_r_shiftReg_28_/7 U9413/4/reg_r_shiftReg_28_/8 U9413/4/46 U9413/4/reg_r_shiftReg_28_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-55.185 19.985 -55.055 20.135)
MU9413/4/reg_r_shiftReg_28_/8 G_DG U9413/4/42 U9413/4/reg_r_shiftReg_28_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-54.705 19.985 -54.575 20.135)
MU9413/4/reg_r_shiftReg_28_/9 U9413/4/reg_r_shiftReg_28_/9 U9413/4/46 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-53.615 19.985 -53.485 20.135)
MU9413/4/reg_r_shiftReg_28_/10 U9413/4/reg_r_shiftReg_28_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_28_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-53.105 19.985 -52.975 20.135)
MU9413/4/reg_r_shiftReg_28_/11 U9413/4/49 U9413/4/42 U9413/4/reg_r_shiftReg_28_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-52.685 19.985 -52.555 20.135)
MU9413/4/reg_r_shiftReg_28_/12 U9413/4/50 U9413/4/49 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-51.595 19.985 -51.465 20.135)
MU9413/4/reg_r_shiftReg_28_/13 U9413/4/51 U9413/4/41 U9413/4/49 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-50.235 19.985 -50.105 20.135)
MU9413/4/reg_r_shiftReg_28_/14 U9413/4/reg_r_shiftReg_28_/14 U9413/4/CLB U9413/4/51 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-49.655 19.985 -49.525 20.135)
MU9413/4/reg_r_shiftReg_28_/15 G_DG U9413/4/50 U9413/4/reg_r_shiftReg_28_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-49.345 19.985 -49.215 20.135)
MU9413/4/reg_r_shiftReg_28_/16 wrData[27] U9413/4/51 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-48.255 19.985 -48.125 20.135)
MU9413/4/reg_r_shiftReg_28_/17 U9413/4/reg_r_shiftReg_28_/QB U9413/4/50 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-47.165 19.985 -47.035 20.135)
MU9413/4/reg_r_shiftReg_30_/1 G_DG U9413/4/CLK U9413/4/28 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-74.635 19.985 -74.505 20.135)
MU9413/4/reg_r_shiftReg_30_/2 U9413/4/29 U9413/4/28 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-74.055 19.985 -73.925 20.135)
MU9413/4/reg_r_shiftReg_30_/3 U9413/4/reg_r_shiftReg_30_/4 U9413/4/ix409/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-72.965 19.985 -72.835 20.135)
MU9413/4/reg_r_shiftReg_30_/4 U9413/4/32 U9413/4/28 U9413/4/reg_r_shiftReg_30_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-72.45 19.985 -72.32 20.135)
MU9413/4/reg_r_shiftReg_30_/5 U9413/4/33 U9413/4/32 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-71.36 19.985 -71.23 20.135)
MU9413/4/reg_r_shiftReg_30_/6 U9413/4/reg_r_shiftReg_30_/7 U9413/4/CLB U9413/4/32 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-69.99 19.985 -69.86 20.135)
MU9413/4/reg_r_shiftReg_30_/7 U9413/4/reg_r_shiftReg_30_/8 U9413/4/33 U9413/4/reg_r_shiftReg_30_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-69.51 19.985 -69.38 20.135)
MU9413/4/reg_r_shiftReg_30_/8 G_DG U9413/4/29 U9413/4/reg_r_shiftReg_30_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-69.03 19.985 -68.9 20.135)
MU9413/4/reg_r_shiftReg_30_/9 U9413/4/reg_r_shiftReg_30_/9 U9413/4/33 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-67.94 19.985 -67.81 20.135)
MU9413/4/reg_r_shiftReg_30_/10 U9413/4/reg_r_shiftReg_30_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_30_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-67.43 19.985 -67.3 20.135)
MU9413/4/reg_r_shiftReg_30_/11 U9413/4/36 U9413/4/29 U9413/4/reg_r_shiftReg_30_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-67.01 19.985 -66.88 20.135)
MU9413/4/reg_r_shiftReg_30_/12 U9413/4/37 U9413/4/36 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-65.92 19.985 -65.79 20.135)
MU9413/4/reg_r_shiftReg_30_/13 U9413/4/38 U9413/4/28 U9413/4/36 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-64.56 19.985 -64.43 20.135)
MU9413/4/reg_r_shiftReg_30_/14 U9413/4/reg_r_shiftReg_30_/14 U9413/4/CLB U9413/4/38 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-63.98 19.985 -63.85 20.135)
MU9413/4/reg_r_shiftReg_30_/15 G_DG U9413/4/37 U9413/4/reg_r_shiftReg_30_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-63.67 19.985 -63.54 20.135)
MU9413/4/reg_r_shiftReg_30_/16 wrData[29] U9413/4/38 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-62.58 19.985 -62.45 20.135)
MU9413/4/reg_r_shiftReg_30_/17 U9413/4/reg_r_shiftReg_30_/QB U9413/4/37 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-61.49 19.985 -61.36 20.135)
MU9413/4/ix409/1 U9413/4/ix409/1 U9413/reg_r_shiftReg_47_\Cross G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-76.395 19.985 -76.265 20.135)
MU9413/4/ix409/2 U9413/4/ix409/OUT U9413/3/ix2027/OUT U9413/4/ix409/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-75.815 19.985 -75.685 20.135)
MU9413/4/reg_r_shiftReg_46_/1 G_DG U9413/4/CLK U9413/4/12 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-90.72 19.985 -90.59 20.135)
MU9413/4/reg_r_shiftReg_46_/2 U9413/4/13 U9413/4/12 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-90.14 19.985 -90.01 20.135)
MU9413/4/reg_r_shiftReg_46_/3 U9413/4/reg_r_shiftReg_46_/4 U9413/4/ix1836/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-89.05 19.985 -88.92 20.135)
MU9413/4/reg_r_shiftReg_46_/4 U9413/4/16 U9413/4/12 U9413/4/reg_r_shiftReg_46_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-88.535 19.985 -88.405 20.135)
MU9413/4/reg_r_shiftReg_46_/5 U9413/4/17 U9413/4/16 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-87.445 19.985 -87.315 20.135)
MU9413/4/reg_r_shiftReg_46_/6 U9413/4/reg_r_shiftReg_46_/7 U9413/4/CLB U9413/4/16 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-86.075 19.985 -85.945 20.135)
MU9413/4/reg_r_shiftReg_46_/7 U9413/4/reg_r_shiftReg_46_/8 U9413/4/17 U9413/4/reg_r_shiftReg_46_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-85.595 19.985 -85.465 20.135)
MU9413/4/reg_r_shiftReg_46_/8 G_DG U9413/4/13 U9413/4/reg_r_shiftReg_46_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-85.115 19.985 -84.985 20.135)
MU9413/4/reg_r_shiftReg_46_/9 U9413/4/reg_r_shiftReg_46_/9 U9413/4/17 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-84.025 19.985 -83.895 20.135)
MU9413/4/reg_r_shiftReg_46_/10 U9413/4/reg_r_shiftReg_46_/10 U9413/4/CLB U9413/4/reg_r_shiftReg_46_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-83.515 19.985 -83.385 20.135)
MU9413/4/reg_r_shiftReg_46_/11 U9413/4/20 U9413/4/13 U9413/4/reg_r_shiftReg_46_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-83.095 19.985 -82.965 20.135)
MU9413/4/reg_r_shiftReg_46_/12 U9413/4/21 U9413/4/20 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-82.005 19.985 -81.875 20.135)
MU9413/4/reg_r_shiftReg_46_/13 U9413/4/22 U9413/4/12 U9413/4/20 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-80.645 19.985 -80.515 20.135)
MU9413/4/reg_r_shiftReg_46_/14 U9413/4/reg_r_shiftReg_46_/14 U9413/4/CLB U9413/4/22 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-80.065 19.985 -79.935 20.135)
MU9413/4/reg_r_shiftReg_46_/15 G_DG U9413/4/21 U9413/4/reg_r_shiftReg_46_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-79.755 19.985 -79.625 20.135)
MU9413/4/reg_r_shiftReg_46_/16 cmd[1] U9413/4/22 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-78.665 19.985 -78.535 20.135)
MU9413/4/reg_r_shiftReg_46_/17 U9413/4/reg_r_shiftReg_46_/QB U9413/4/21 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-77.575 19.985 -77.445 20.135)
MU9413/4/ix1836/1 G_DG U9413/SEL U9413/4/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-94.8 19.985 -94.67 20.135)
MU9413/4/ix1836/2 U9413/4/ix1836/3 U9413/4/5 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-94.22 19.985 -94.09 20.135)
MU9413/4/ix1836/3 U9413/4/7 cmd[1] U9413/4/ix1836/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-93.64 19.985 -93.51 20.135)
MU9413/4/ix1836/4 U9413/4/ix1836/5 cmd[0] U9413/4/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-93.06 19.985 -92.93 20.135)
MU9413/4/ix1836/5 G_DG U9413/SEL U9413/4/ix1836/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-92.48 19.985 -92.35 20.135)
MU9413/4/ix1836/6 U9413/4/ix1836/OUT U9413/4/7 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-91.9 19.985 -91.77 20.135)
MU9413/5/1 G_DS CLK U9413/5/2 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-98.32 13.22 -98.19 13.52)
MU9413/5/2 U9413/5/CLK U9413/5/2 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-97.74 13.22 -97.61 13.52)
MU9413/5/3 G_DS CLK U9413/5/3 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-96.56 13.22 -96.43 13.52)
MU9413/5/4 U9413/5/CLK U9413/5/3 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-95.98 13.22 -95.85 13.52)
MU9413/5/5 G_DS CLK U9413/5/4 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-94.8 13.22 -94.67 13.52)
MU9413/5/6 U9413/5/CLK U9413/5/4 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-94.22 13.22 -94.09 13.52)
MU9413/5/7 G_DS U9413/SEL U9413/5/6 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-93.04 13.005 -92.91 13.305)
MU9413/5/8 U9413/5/7 U9413/5/6 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-92.46 13.005 -92.33 13.525)
MU9413/5/9 U9413/5/8 cmd[2] U9413/5/7 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-91.88 13.005 -91.75 13.525)
MU9413/5/10 U9413/5/10 cmd[3] U9413/5/8 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-91.3 13.005 -91.17 13.525)
MU9413/5/11 G_DS U9413/SEL U9413/5/10 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-90.72 13.005 -90.59 13.525)
MU9413/5/12 U9413/5/ix1856/OUT U9413/5/8 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-90.14 13.22 -90.01 13.52)
MU9413/5/13 G_DS U9413/5/ix1876/SEL U9413/5/14 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-88.96 13.005 -88.83 13.305)
MU9413/5/14 U9413/5/15 U9413/5/14 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-88.38 13.005 -88.25 13.525)
MU9413/5/15 U9413/5/16 cmd[4] U9413/5/15 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-87.8 13.005 -87.67 13.525)
MU9413/5/16 U9413/5/18 cmd[5] U9413/5/16 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-87.22 13.005 -87.09 13.525)
MU9413/5/17 G_DS U9413/5/ix1876/SEL U9413/5/18 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-86.64 13.005 -86.51 13.525)
MU9413/5/18 U9413/5/ix1876/OUT U9413/5/16 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-86.06 13.22 -85.93 13.52)
MU9413/5/19 G_DS U9413/5/CLK U9413/5/21 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-84.88 13.22 -84.75 13.52)
MU9413/5/20 U9413/5/22 U9413/5/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-84.3 13.22 -84.17 13.52)
MU9413/5/21 U9413/5/23 U9413/5/ix1876/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-83.21 13.22 -83.08 13.61)
MU9413/5/22 U9413/5/25 U9413/5/22 U9413/5/23 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-82.695 13.22 -82.565 13.61)
MU9413/5/23 U9413/5/26 U9413/5/25 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-81.605 13.22 -81.475 13.52)
MU9413/5/24 U9413/5/27 U9413/5/21 U9413/5/25 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-80.515 13.22 -80.385 13.61)
MU9413/5/25 G_DS U9413/5/CLB U9413/5/27 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-79.895 13.22 -79.765 13.61)
MU9413/5/26 U9413/5/27 U9413/5/26 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-79.275 13.22 -79.145 13.61)
MU9413/5/27 U9413/5/28 U9413/5/26 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-78.185 13.22 -78.055 13.61)
MU9413/5/28 U9413/5/29 U9413/5/21 U9413/5/28 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-77.875 13.22 -77.745 13.61)
MU9413/5/29 U9413/5/30 U9413/5/29 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-76.165 13.22 -76.035 13.52)
MU9413/5/30 U9413/5/31 U9413/5/22 U9413/5/29 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-75.075 13.22 -74.945 13.61)
MU9413/5/31 G_DS U9413/5/CLB U9413/5/31 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-74.495 13.22 -74.365 13.61)
MU9413/5/32 U9413/5/31 U9413/5/30 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-73.915 13.22 -73.785 13.52)
MU9413/5/33 cmd[5] U9413/5/31 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-72.825 13.22 -72.695 13.52)
MU9413/5/34 U9413/5/reg_r_shiftReg_50_/QB U9413/5/30 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-71.735 13.22 -71.605 13.52)
MU9413/5/35 G_DS U9413/5/ix1876/SEL U9413/5/35 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-70.555 13.005 -70.425 13.305)
MU9413/5/36 U9413/5/36 U9413/5/35 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-69.975 13.005 -69.845 13.525)
MU9413/5/37 U9413/5/37 cmd[5] U9413/5/36 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-69.395 13.005 -69.265 13.525)
MU9413/5/38 U9413/5/39 cmd[6] U9413/5/37 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-68.815 13.005 -68.685 13.525)
MU9413/5/39 G_DS U9413/5/ix1876/SEL U9413/5/39 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-68.235 13.005 -68.105 13.525)
MU9413/5/40 U9413/5/ix1886/OUT U9413/5/37 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-67.655 13.22 -67.525 13.52)
MU9413/5/41 G_DS U9413/5/CLK U9413/5/42 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-66.475 13.22 -66.345 13.52)
MU9413/5/42 U9413/5/43 U9413/5/42 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-65.895 13.22 -65.765 13.52)
MU9413/5/43 U9413/5/44 U9413/5/ix1886/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-64.805 13.22 -64.675 13.61)
MU9413/5/44 U9413/5/46 U9413/5/43 U9413/5/44 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-64.29 13.22 -64.16 13.61)
MU9413/5/45 U9413/5/47 U9413/5/46 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-63.2 13.22 -63.07 13.52)
MU9413/5/46 U9413/5/48 U9413/5/42 U9413/5/46 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-62.11 13.22 -61.98 13.61)
MU9413/5/47 G_DS U9413/5/CLB U9413/5/48 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-61.49 13.22 -61.36 13.61)
MU9413/5/48 U9413/5/48 U9413/5/47 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-60.87 13.22 -60.74 13.61)
MU9413/5/49 U9413/5/49 U9413/5/47 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-59.78 13.22 -59.65 13.61)
MU9413/5/50 U9413/5/50 U9413/5/42 U9413/5/49 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-59.47 13.22 -59.34 13.61)
MU9413/5/51 U9413/5/51 U9413/5/50 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-57.76 13.22 -57.63 13.52)
MU9413/5/52 U9413/5/52 U9413/5/43 U9413/5/50 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-56.67 13.22 -56.54 13.61)
MU9413/5/53 G_DS U9413/5/CLB U9413/5/52 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-56.09 13.22 -55.96 13.61)
MU9413/5/54 U9413/5/52 U9413/5/51 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-55.51 13.22 -55.38 13.52)
MU9413/5/55 cmd[6] U9413/5/52 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-54.42 13.22 -54.29 13.52)
MU9413/5/56 U9413/5/reg_r_shiftReg_51_/QB U9413/5/51 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-53.33 13.22 -53.2 13.52)
MU9413/5/57 G_DS U9413/5/ix1916/SEL U9413/5/56 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-52.15 13.005 -52.02 13.305)
MU9413/5/58 U9413/5/57 U9413/5/56 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-51.57 13.005 -51.44 13.525)
MU9413/5/59 U9413/5/58 cmd[6] U9413/5/57 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-50.99 13.005 -50.86 13.525)
MU9413/5/60 U9413/5/60 readL U9413/5/58 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-50.41 13.005 -50.28 13.525)
MU9413/5/61 G_DS U9413/5/ix1916/SEL U9413/5/60 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-49.83 13.005 -49.7 13.525)
MU9413/5/62 U9413/5/ix1916/OUT U9413/5/58 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-49.25 13.22 -49.12 13.52)
MU9413/5/63 G_DS U9413/5/ix1876/SEL U9413/5/64 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-48.07 13.005 -47.94 13.305)
MU9413/5/64 U9413/5/65 U9413/5/64 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-47.49 13.005 -47.36 13.525)
MU9413/5/65 U9413/5/66 cmd[6] U9413/5/65 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-46.91 13.005 -46.78 13.525)
MU9413/5/66 U9413/5/68 U9413/5/ix1896/B U9413/5/66 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-46.33 13.005 -46.2 13.525)
MU9413/5/67 G_DS U9413/5/ix1876/SEL U9413/5/68 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-45.75 13.005 -45.62 13.525)
MU9413/5/68 U9413/5/ix1896/OUT U9413/5/66 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-45.17 13.22 -45.04 13.52)
MU9413/5/69 U9413/5/71 exec G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-43.99 13.005 -43.86 13.525)
MU9413/5/70 U9413/5/73 U9413/5/ix489/B U9413/5/71 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.17e-013 pd=9.7e-007 ps=9.7e-007 nrd=0.432692 nrs=0.432692  $(-43.41 13.005 -43.28 13.525)
MU9413/5/71 U9413/5/ix1916/SEL U9413/5/ix489/C U9413/5/73 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-42.83 13.005 -42.7 13.525)
MU9413/5/72 G_DS U9413/5/CLK U9413/5/77 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-41.65 13.22 -41.52 13.52)
MU9413/5/73 U9413/5/78 U9413/5/77 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-41.07 13.22 -40.94 13.52)
MU9413/5/74 U9413/5/79 U9413/5/ix1896/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-39.98 13.22 -39.85 13.61)
MU9413/5/75 U9413/5/81 U9413/5/78 U9413/5/79 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-39.465 13.22 -39.335 13.61)
MU9413/5/76 U9413/5/82 U9413/5/81 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-38.375 13.22 -38.245 13.52)
MU9413/5/77 U9413/5/83 U9413/5/77 U9413/5/81 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-37.285 13.22 -37.155 13.61)
MU9413/5/78 G_DS U9413/5/CLB U9413/5/83 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-36.665 13.22 -36.535 13.61)
MU9413/5/79 U9413/5/83 U9413/5/82 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-36.045 13.22 -35.915 13.61)
MU9413/5/80 U9413/5/84 U9413/5/82 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-34.955 13.22 -34.825 13.61)
MU9413/5/81 U9413/5/85 U9413/5/77 U9413/5/84 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-34.645 13.22 -34.515 13.61)
MU9413/5/82 U9413/5/86 U9413/5/85 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-32.935 13.22 -32.805 13.52)
MU9413/5/83 U9413/5/87 U9413/5/78 U9413/5/85 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-31.845 13.22 -31.715 13.61)
MU9413/5/84 G_DS U9413/5/CLB U9413/5/87 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-31.265 13.22 -31.135 13.61)
MU9413/5/85 U9413/5/87 U9413/5/86 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-30.685 13.22 -30.555 13.52)
MU9413/5/86 U9413/5/ix1896/B U9413/5/87 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-29.595 13.22 -29.465 13.52)
MU9413/5/87 U9413/5/ix489/C U9413/5/86 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-28.505 13.22 -28.375 13.52)
MU9413/5/88 G_DS U9413/4/ix2270/A U9413/5/91 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-27.325 13.22 -27.195 13.52)
MU9413/5/89 U9413/5/ix1876/SEL U9413/5/91 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-26.745 13.22 -26.615 13.52)
MU9413/5/90 U9413/4/ix2270/A exec G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-25.565 13.22 -25.435 13.48)
MU9413/5/91 G_DS U9413/5/C U9413/4/ix2270/A G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(-24.985 13.22 -24.855 13.48)
MU9413/5/92 G_DS U9413/5/CLK U9413/5/96 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-23.805 13.22 -23.675 13.52)
MU9413/5/93 U9413/5/97 U9413/5/96 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-23.225 13.22 -23.095 13.52)
MU9413/5/94 U9413/5/98 U9413/5/ix25/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-22.135 13.22 -22.005 13.61)
MU9413/5/95 U9413/5/100 U9413/5/97 U9413/5/98 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-21.62 13.22 -21.49 13.61)
MU9413/5/96 U9413/5/101 U9413/5/100 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-20.53 13.22 -20.4 13.52)
MU9413/5/97 U9413/5/102 U9413/5/96 U9413/5/100 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-19.44 13.22 -19.31 13.61)
MU9413/5/98 G_DS U9413/5/CLB U9413/5/102 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-18.82 13.22 -18.69 13.61)
MU9413/5/99 U9413/5/102 U9413/5/101 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-18.2 13.22 -18.07 13.61)
MU9413/5/100 U9413/5/103 U9413/5/101 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-17.11 13.22 -16.98 13.61)
MU9413/5/101 U9413/5/104 U9413/5/96 U9413/5/103 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-16.8 13.22 -16.67 13.61)
MU9413/5/102 U9413/5/105 U9413/5/104 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-15.09 13.22 -14.96 13.52)
MU9413/5/103 U9413/5/106 U9413/5/97 U9413/5/104 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-14 13.22 -13.87 13.61)
MU9413/5/104 G_DS U9413/5/CLB U9413/5/106 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-13.42 13.22 -13.29 13.61)
MU9413/5/105 U9413/5/106 U9413/5/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-12.84 13.22 -12.71 13.52)
MU9413/5/106 U9413/5/C U9413/5/106 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-11.75 13.22 -11.62 13.52)
MU9413/5/107 U9413/5/ix489/B U9413/5/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-10.66 13.22 -10.53 13.52)
MU9413/5/108 U9413/5/109 U9413/5/ix1896/B G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-9.48 13.005 -9.35 13.525)
MU9413/5/109 U9413/5/111 U9413/5/ix2004/OUT U9413/5/109 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.17e-013 pd=9.7e-007 ps=9.7e-007 nrd=0.432692 nrs=0.432692  $(-8.9 13.005 -8.77 13.525)
MU9413/5/110 U9413/3/ix2292/A U9413/5/ix489/B U9413/5/111 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-8.32 13.005 -8.19 13.525)
MU9413/5/111 U9413/5/ix2004/OUT ack G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-7.14 13.22 -7.01 13.52)
MU9413/5/112 G_DS U9413/QB U9413/5/118 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-5.96 13.005 -5.83 13.305)
MU9413/5/113 U9413/5/119 U9413/5/118 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-5.38 13.005 -5.25 13.525)
MU9413/5/114 U9413/5/120 U9413/4/ix2251/A U9413/5/119 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-4.8 13.005 -4.67 13.525)
MU9413/5/115 U9413/5/122 U9413/5/ix2004/OUT U9413/5/120 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-4.22 13.005 -4.09 13.525)
MU9413/5/116 G_DS U9413/QB U9413/5/122 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-3.64 13.005 -3.51 13.525)
MU9413/5/117 U9413/5/ix25/OUT U9413/5/120 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-3.06 13.22 -2.93 13.52)
MU9413/5/118 U9413/5/ix2272/A exec G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(0.47 13.22 0.6 13.48)
MU9413/5/119 G_DS U9413/5/C U9413/5/ix2272/A G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(1.05 13.22 1.18 13.48)
MU9413/5/120 U9413/4/ix2276/A U9413/5/ix2198/OUT G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(2.23 13.22 2.36 13.48)
MU9413/5/121 G_DS U9413/5/ix39/B U9413/4/ix2276/A G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=1.365e-013 pd=1.53e-006 ps=8.4e-007 nrd=2.01923 nrs=1.15385  $(2.81 13.22 2.94 13.48)
MU9413/5/122 G_DS U9413/5/CLK U9413/5/131 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(3.99 13.22 4.12 13.52)
MU9413/5/123 U9413/5/132 U9413/5/131 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(4.57 13.22 4.7 13.52)
MU9413/5/124 U9413/5/133 U9413/5/ix25/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(5.66 13.22 5.79 13.61)
MU9413/5/125 U9413/5/135 U9413/5/132 U9413/5/133 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(6.175 13.22 6.305 13.61)
MU9413/5/126 U9413/5/136 U9413/5/135 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(7.265 13.22 7.395 13.52)
MU9413/5/127 U9413/5/137 U9413/5/131 U9413/5/135 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(8.355 13.22 8.485 13.61)
MU9413/5/128 G_DS U9413/5/CLB U9413/5/137 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(8.975 13.22 9.105 13.61)
MU9413/5/129 U9413/5/137 U9413/5/136 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(9.595 13.22 9.725 13.61)
MU9413/5/130 U9413/5/138 U9413/5/136 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(10.685 13.22 10.815 13.61)
MU9413/5/131 U9413/5/139 U9413/5/131 U9413/5/138 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(10.995 13.22 11.125 13.61)
MU9413/5/132 U9413/5/140 U9413/5/139 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(12.705 13.22 12.835 13.52)
MU9413/5/133 U9413/5/141 U9413/5/132 U9413/5/139 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(13.795 13.22 13.925 13.61)
MU9413/5/134 G_DS U9413/5/CLB U9413/5/141 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(14.375 13.22 14.505 13.61)
MU9413/5/135 U9413/5/141 U9413/5/140 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(14.955 13.22 15.085 13.52)
MU9413/5/136 U9413/5/ix39/B U9413/5/141 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(16.045 13.22 16.175 13.52)
MU9413/5/137 U9413/QB U9413/5/140 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(17.135 13.22 17.265 13.52)
MU9413/5/138 G_DS U9413/5/ix2272/A U9413/5/144 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(18.315 13.22 18.445 13.52)
MU9413/5/139 U9413/6/SEL U9413/5/144 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(18.895 13.22 19.025 13.52)
MU9413/5/140 G_DS U9413/5/ix2272/A U9413/5/147 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(20.075 13.22 20.205 13.52)
MU9413/5/141 U9413/SEL U9413/5/147 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(20.655 13.22 20.785 13.52)
MU9413/5/142 G_DS U9413/5/CLK U9413/5/149 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(21.835 13.22 21.965 13.52)
MU9413/5/143 U9413/5/150 U9413/5/149 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(22.415 13.22 22.545 13.52)
MU9413/5/144 U9413/5/151 U9413/5/reg_r_shiftReg_0_/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(23.505 13.22 23.635 13.61)
MU9413/5/145 U9413/5/153 U9413/5/150 U9413/5/151 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(24.02 13.22 24.15 13.61)
MU9413/5/146 U9413/5/154 U9413/5/153 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(25.11 13.22 25.24 13.52)
MU9413/5/147 U9413/5/155 U9413/5/149 U9413/5/153 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(26.2 13.22 26.33 13.61)
MU9413/5/148 G_DS U9413/5/CLB U9413/5/155 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(26.82 13.22 26.95 13.61)
MU9413/5/149 U9413/5/155 U9413/5/154 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(27.44 13.22 27.57 13.61)
MU9413/5/150 U9413/5/156 U9413/5/154 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(28.53 13.22 28.66 13.61)
MU9413/5/151 U9413/5/157 U9413/5/149 U9413/5/156 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(28.84 13.22 28.97 13.61)
MU9413/5/152 U9413/5/158 U9413/5/157 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(30.55 13.22 30.68 13.52)
MU9413/5/153 U9413/5/159 U9413/5/150 U9413/5/157 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(31.64 13.22 31.77 13.61)
MU9413/5/154 G_DS U9413/5/CLB U9413/5/159 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(32.22 13.22 32.35 13.61)
MU9413/5/155 U9413/5/159 U9413/5/158 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(32.8 13.22 32.93 13.52)
MU9413/5/156 U9413/4/ix2251/A U9413/5/159 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(33.89 13.22 34.02 13.52)
MU9413/5/157 U9413/5/reg_r_shiftReg_0_/QB U9413/5/158 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(34.98 13.22 35.11 13.52)
MU9413/5/158 G_DS U9413/5/CLK U9413/5/162 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(36.16 13.22 36.29 13.52)
MU9413/5/159 U9413/5/163 U9413/5/162 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(36.74 13.22 36.87 13.52)
MU9413/5/160 U9413/5/164 U9413/4/ix229/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(37.83 13.22 37.96 13.61)
MU9413/5/161 U9413/5/166 U9413/5/163 U9413/5/164 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(38.345 13.22 38.475 13.61)
MU9413/5/162 U9413/5/167 U9413/5/166 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(39.435 13.22 39.565 13.52)
MU9413/5/163 U9413/5/168 U9413/5/162 U9413/5/166 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(40.525 13.22 40.655 13.61)
MU9413/5/164 G_DS U9413/5/CLB U9413/5/168 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(41.145 13.22 41.275 13.61)
MU9413/5/165 U9413/5/168 U9413/5/167 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(41.765 13.22 41.895 13.61)
MU9413/5/166 U9413/5/169 U9413/5/167 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(42.855 13.22 42.985 13.61)
MU9413/5/167 U9413/5/170 U9413/5/162 U9413/5/169 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(43.165 13.22 43.295 13.61)
MU9413/5/168 U9413/5/171 U9413/5/170 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(44.875 13.22 45.005 13.52)
MU9413/5/169 U9413/5/172 U9413/5/163 U9413/5/170 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(45.965 13.22 46.095 13.61)
MU9413/5/170 G_DS U9413/5/CLB U9413/5/172 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(46.545 13.22 46.675 13.61)
MU9413/5/171 U9413/5/172 U9413/5/171 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(47.125 13.22 47.255 13.52)
MU9413/5/172 wrData[14] U9413/5/172 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(48.215 13.22 48.345 13.52)
MU9413/5/173 U9413/5/reg_r_shiftReg_15_/QB U9413/5/171 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(49.305 13.22 49.435 13.52)
MU9413/5/174 G_DS U9413/SEL U9413/5/176 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(50.485 13.005 50.615 13.305)
MU9413/5/175 U9413/5/177 U9413/5/176 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(51.065 13.005 51.195 13.525)
MU9413/5/176 U9413/5/178 addr[11] U9413/5/177 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(51.645 13.005 51.775 13.525)
MU9413/5/177 U9413/5/180 cmd[0] U9413/5/178 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(52.225 13.005 52.355 13.525)
MU9413/5/178 G_DS U9413/SEL U9413/5/180 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(52.805 13.005 52.935 13.525)
MU9413/5/179 U9413/5/ix1826/OUT U9413/5/178 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(53.385 13.22 53.515 13.52)
MU9413/5/180 G_DS U9413/5/CLK U9413/5/183 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(54.565 13.22 54.695 13.52)
MU9413/5/181 U9413/5/184 U9413/5/183 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(55.145 13.22 55.275 13.52)
MU9413/5/182 U9413/5/185 U9413/4/ix205/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(56.235 13.22 56.365 13.61)
MU9413/5/183 U9413/5/187 U9413/5/184 U9413/5/185 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(56.75 13.22 56.88 13.61)
MU9413/5/184 U9413/5/188 U9413/5/187 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(57.84 13.22 57.97 13.52)
MU9413/5/185 U9413/5/189 U9413/5/183 U9413/5/187 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(58.93 13.22 59.06 13.61)
MU9413/5/186 G_DS U9413/5/CLB U9413/5/189 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(59.55 13.22 59.68 13.61)
MU9413/5/187 U9413/5/189 U9413/5/188 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(60.17 13.22 60.3 13.61)
MU9413/5/188 U9413/5/190 U9413/5/188 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(61.26 13.22 61.39 13.61)
MU9413/5/189 U9413/5/191 U9413/5/183 U9413/5/190 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(61.57 13.22 61.7 13.61)
MU9413/5/190 U9413/5/192 U9413/5/191 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(63.28 13.22 63.41 13.52)
MU9413/5/191 U9413/5/193 U9413/5/184 U9413/5/191 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(64.37 13.22 64.5 13.61)
MU9413/5/192 G_DS U9413/5/CLB U9413/5/193 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(64.95 13.22 65.08 13.61)
MU9413/5/193 U9413/5/193 U9413/5/192 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(65.53 13.22 65.66 13.52)
MU9413/5/194 wrData[12] U9413/5/193 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(66.62 13.22 66.75 13.52)
MU9413/5/195 U9413/5/reg_r_shiftReg_13_/QB U9413/5/192 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(67.71 13.22 67.84 13.52)
MU9413/5/196 G_DS U9413/5/CLK U9413/5/196 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(68.89 13.22 69.02 13.52)
MU9413/5/197 U9413/5/197 U9413/5/196 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(69.47 13.22 69.6 13.52)
MU9413/5/198 U9413/5/198 U9413/4/ix145/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(70.56 13.22 70.69 13.61)
MU9413/5/199 U9413/5/200 U9413/5/197 U9413/5/198 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(71.075 13.22 71.205 13.61)
MU9413/5/200 U9413/5/201 U9413/5/200 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(72.165 13.22 72.295 13.52)
MU9413/5/201 U9413/5/202 U9413/5/196 U9413/5/200 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(73.255 13.22 73.385 13.61)
MU9413/5/202 G_DS U9413/5/CLB U9413/5/202 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(73.875 13.22 74.005 13.61)
MU9413/5/203 U9413/5/202 U9413/5/201 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(74.495 13.22 74.625 13.61)
MU9413/5/204 U9413/5/203 U9413/5/201 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(75.585 13.22 75.715 13.61)
MU9413/5/205 U9413/5/204 U9413/5/196 U9413/5/203 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(75.895 13.22 76.025 13.61)
MU9413/5/206 U9413/5/205 U9413/5/204 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(77.605 13.22 77.735 13.52)
MU9413/5/207 U9413/5/206 U9413/5/197 U9413/5/204 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(78.695 13.22 78.825 13.61)
MU9413/5/208 G_DS U9413/5/CLB U9413/5/206 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(79.275 13.22 79.405 13.61)
MU9413/5/209 U9413/5/206 U9413/5/205 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(79.855 13.22 79.985 13.52)
MU9413/5/210 wrData[7] U9413/5/206 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(80.945 13.22 81.075 13.52)
MU9413/5/211 U9413/5/reg_r_shiftReg_8_/QB U9413/5/205 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(82.035 13.22 82.165 13.52)
MU9413/5/212 G_DS U9413/5/CLK U9413/5/209 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(83.215 13.22 83.345 13.52)
MU9413/5/213 U9413/5/210 U9413/5/209 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(83.795 13.22 83.925 13.52)
MU9413/5/214 U9413/5/211 U9413/5/reg_r_shiftReg_35_/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(84.885 13.22 85.015 13.61)
MU9413/5/215 U9413/5/213 U9413/5/210 U9413/5/211 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(85.4 13.22 85.53 13.61)
MU9413/5/216 U9413/5/214 U9413/5/213 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(86.49 13.22 86.62 13.52)
MU9413/5/217 U9413/5/215 U9413/5/209 U9413/5/213 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(87.58 13.22 87.71 13.61)
MU9413/5/218 G_DS U9413/5/CLB U9413/5/215 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(88.2 13.22 88.33 13.61)
MU9413/5/219 U9413/5/215 U9413/5/214 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(88.82 13.22 88.95 13.61)
MU9413/5/220 U9413/5/216 U9413/5/214 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(89.91 13.22 90.04 13.61)
MU9413/5/221 U9413/5/217 U9413/5/209 U9413/5/216 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(90.22 13.22 90.35 13.61)
MU9413/5/222 U9413/5/218 U9413/5/217 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(91.93 13.22 92.06 13.52)
MU9413/5/223 U9413/5/219 U9413/5/210 U9413/5/217 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(93.02 13.22 93.15 13.61)
MU9413/5/224 G_DS U9413/5/CLB U9413/5/219 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(93.6 13.22 93.73 13.61)
MU9413/5/225 U9413/5/219 U9413/5/218 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(94.18 13.22 94.31 13.52)
MU9413/5/226 addr[2] U9413/5/219 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(95.27 13.22 95.4 13.52)
MU9413/5/227 U9413/5/reg_r_shiftReg_35_/QB U9413/5/218 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(96.36 13.22 96.49 13.52)
MU9413/5/228 U9413/5/222 ack G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(97.54 13.005 97.67 13.525)
MU9413/5/229 U9413/D U9413/6/SEL U9413/5/222 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(98.12 13.005 98.25 13.525)
MU9413/5/230 G_DS U9413/5/CLK U9413/5/226 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(99.3 13.22 99.43 13.52)
MU9413/5/231 U9413/5/227 U9413/5/226 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(99.88 13.22 100.01 13.52)
MU9413/5/232 U9413/5/228 U9413/ix1786\Cross G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(100.97 13.22 101.1 13.61)
MU9413/5/233 U9413/5/230 U9413/5/227 U9413/5/228 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(101.485 13.22 101.615 13.61)
MU9413/5/234 U9413/5/231 U9413/5/230 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(102.575 13.22 102.705 13.52)
MU9413/5/235 U9413/5/232 U9413/5/226 U9413/5/230 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(103.665 13.22 103.795 13.61)
MU9413/5/236 G_DS U9413/5/CLB U9413/5/232 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(104.285 13.22 104.415 13.61)
MU9413/5/237 U9413/5/232 U9413/5/231 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(104.905 13.22 105.035 13.61)
MU9413/5/238 U9413/5/233 U9413/5/231 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(105.995 13.22 106.125 13.61)
MU9413/5/239 U9413/5/234 U9413/5/226 U9413/5/233 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(106.305 13.22 106.435 13.61)
MU9413/5/240 U9413/5/235 U9413/5/234 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(108.015 13.22 108.145 13.52)
MU9413/5/241 U9413/5/236 U9413/5/227 U9413/5/234 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(109.105 13.22 109.235 13.61)
MU9413/5/242 G_DS U9413/5/CLB U9413/5/236 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(109.685 13.22 109.815 13.61)
MU9413/5/243 U9413/5/236 U9413/5/235 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(110.265 13.22 110.395 13.52)
MU9413/5/244 wrData[2] U9413/5/236 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(111.355 13.22 111.485 13.52)
MU9413/5/245 U9413/5/reg_r_shiftReg_3_/QB U9413/5/235 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(112.445 13.22 112.575 13.52)
MU9413/5/246 G_DS U9413/5/CLK U9413/5/239 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(113.625 13.22 113.755 13.52)
MU9413/5/247 U9413/5/240 U9413/5/239 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(114.205 13.22 114.335 13.52)
MU9413/5/248 U9413/5/241 U9413/5/ix1766/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(115.295 13.22 115.425 13.61)
MU9413/5/249 U9413/5/243 U9413/5/240 U9413/5/241 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(115.81 13.22 115.94 13.61)
MU9413/5/250 U9413/5/244 U9413/5/243 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(116.9 13.22 117.03 13.52)
MU9413/5/251 U9413/5/245 U9413/5/239 U9413/5/243 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(117.99 13.22 118.12 13.61)
MU9413/5/252 G_DS U9413/5/CLB U9413/5/245 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(118.61 13.22 118.74 13.61)
MU9413/5/253 U9413/5/245 U9413/5/244 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(119.23 13.22 119.36 13.61)
MU9413/5/254 U9413/5/246 U9413/5/244 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(120.32 13.22 120.45 13.61)
MU9413/5/255 U9413/5/247 U9413/5/239 U9413/5/246 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(120.63 13.22 120.76 13.61)
MU9413/5/256 U9413/5/248 U9413/5/247 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(122.34 13.22 122.47 13.52)
MU9413/5/257 U9413/5/249 U9413/5/240 U9413/5/247 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(123.43 13.22 123.56 13.61)
MU9413/5/258 G_DS U9413/5/CLB U9413/5/249 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(124.01 13.22 124.14 13.61)
MU9413/5/259 U9413/5/249 U9413/5/248 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(124.59 13.22 124.72 13.52)
MU9413/5/260 addr[6] U9413/5/249 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(125.68 13.22 125.81 13.52)
MU9413/5/261 U9413/5/reg_r_shiftReg_39_/QB U9413/5/248 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(126.77 13.22 126.9 13.52)
MU9413/5/262 G_DS U9413/6/SEL U9413/5/253 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(127.95 13.005 128.08 13.305)
MU9413/5/263 U9413/5/254 U9413/5/253 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(128.53 13.005 128.66 13.525)
MU9413/5/264 U9413/5/255 addr[5] U9413/5/254 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(129.11 13.005 129.24 13.525)
MU9413/5/265 U9413/5/257 addr[6] U9413/5/255 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(129.69 13.005 129.82 13.525)
MU9413/5/266 G_DS U9413/6/SEL U9413/5/257 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(130.27 13.005 130.4 13.525)
MU9413/5/267 U9413/5/ix1766/OUT U9413/5/255 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(130.85 13.22 130.98 13.52)
MU9413/5/268 G_DS U9413/SEL U9413/5/260 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(132.03 13.005 132.16 13.305)
MU9413/5/269 U9413/5/261 U9413/5/260 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(132.61 13.005 132.74 13.525)
MU9413/5/270 U9413/5/262 addr[6] U9413/5/261 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(133.19 13.005 133.32 13.525)
MU9413/5/271 U9413/5/263 addr[7] U9413/5/262 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(133.77 13.005 133.9 13.525)
MU9413/5/272 G_DS U9413/SEL U9413/5/263 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(134.35 13.005 134.48 13.525)
MU9413/5/273 U9413/5/DATA U9413/5/262 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(134.93 13.22 135.06 13.52)
MU9413/5/274 G_DS U9413/5/CLK U9413/5/264 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(136.11 13.22 136.24 13.52)
MU9413/5/275 U9413/5/265 U9413/5/264 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(136.69 13.22 136.82 13.52)
MU9413/5/276 U9413/5/266 U9413/5/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(137.78 13.22 137.91 13.61)
MU9413/5/277 U9413/5/267 U9413/5/265 U9413/5/266 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(138.295 13.22 138.425 13.61)
MU9413/5/278 U9413/5/268 U9413/5/267 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(139.385 13.22 139.515 13.52)
MU9413/5/279 U9413/5/269 U9413/5/264 U9413/5/267 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(140.475 13.22 140.605 13.61)
MU9413/5/280 G_DS U9413/5/CLB U9413/5/269 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(141.095 13.22 141.225 13.61)
MU9413/5/281 U9413/5/269 U9413/5/268 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(141.715 13.22 141.845 13.61)
MU9413/5/282 U9413/5/270 U9413/5/268 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(142.805 13.22 142.935 13.61)
MU9413/5/283 U9413/5/271 U9413/5/264 U9413/5/270 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(143.115 13.22 143.245 13.61)
MU9413/5/284 U9413/5/272 U9413/5/271 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(144.825 13.22 144.955 13.52)
MU9413/5/285 U9413/5/273 U9413/5/265 U9413/5/271 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(145.915 13.22 146.045 13.61)
MU9413/5/286 G_DS U9413/5/CLB U9413/5/273 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(146.495 13.22 146.625 13.61)
MU9413/5/287 U9413/5/273 U9413/5/272 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(147.075 13.22 147.205 13.52)
MU9413/5/288 addr[7] U9413/5/273 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(148.165 13.22 148.295 13.52)
MU9413/5/289 U9413/5/reg_r_shiftReg_40_/QB U9413/5/272 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(149.255 13.22 149.385 13.52)
MU9413/5/290 G_DS RST U9413/5/275 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(150.435 13.22 150.565 13.52)
MU9413/5/291 U9413/5/CLB U9413/5/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(151.015 13.22 151.145 13.52)
MU9413/5/292 G_DS RST U9413/5/276 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(152.195 13.22 152.325 13.52)
MU9413/5/293 U9413/5/CLB U9413/5/276 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(152.775 13.22 152.905 13.52)
MU9413/5/294 G_DS RST U9413/5/277 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(153.955 13.22 154.085 13.52)
MU9413/5/295 U9413/5/CLB U9413/5/277 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(154.535 13.22 154.665 13.52)
MU9413/5/right_22/1 G_DG RST U9413/5/275 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(150.435 11.49 150.565 11.64)
MU9413/5/right_22/2 U9413/5/CLB U9413/5/275 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(151.015 11.49 151.145 11.64)
MU9413/5/right_21/1 G_DG RST U9413/5/276 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(152.195 11.49 152.325 11.64)
MU9413/5/right_21/2 U9413/5/CLB U9413/5/276 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(152.775 11.49 152.905 11.64)
MU9413/5/right_20/1 G_DG RST U9413/5/277 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(153.955 11.49 154.085 11.64)
MU9413/5/right_20/2 U9413/5/CLB U9413/5/277 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(154.535 11.49 154.665 11.64)
MU9413/5/left_22/1 G_DG CLK U9413/5/2 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-98.32 11.49 -98.19 11.64)
MU9413/5/left_22/2 U9413/5/CLK U9413/5/2 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-97.74 11.49 -97.61 11.64)
MU9413/5/left_21/1 G_DG CLK U9413/5/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-96.56 11.49 -96.43 11.64)
MU9413/5/left_21/2 U9413/5/CLK U9413/5/3 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-95.98 11.49 -95.85 11.64)
MU9413/5/left_20/1 G_DG CLK U9413/5/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-94.8 11.49 -94.67 11.64)
MU9413/5/left_20/2 U9413/5/CLK U9413/5/4 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-94.22 11.49 -94.09 11.64)
MU9413/5/reg_r_shiftReg_40_/1 G_DG U9413/5/CLK U9413/5/264 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(136.11 11.49 136.24 11.64)
MU9413/5/reg_r_shiftReg_40_/2 U9413/5/265 U9413/5/264 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(136.69 11.49 136.82 11.64)
MU9413/5/reg_r_shiftReg_40_/3 U9413/5/reg_r_shiftReg_40_/4 U9413/5/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(137.78 11.49 137.91 11.64)
MU9413/5/reg_r_shiftReg_40_/4 U9413/5/267 U9413/5/264 U9413/5/reg_r_shiftReg_40_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(138.295 11.49 138.425 11.64)
MU9413/5/reg_r_shiftReg_40_/5 U9413/5/268 U9413/5/267 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(139.385 11.49 139.515 11.64)
MU9413/5/reg_r_shiftReg_40_/6 U9413/5/reg_r_shiftReg_40_/7 U9413/5/CLB U9413/5/267 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(140.755 11.49 140.885 11.64)
MU9413/5/reg_r_shiftReg_40_/7 U9413/5/reg_r_shiftReg_40_/8 U9413/5/268 U9413/5/reg_r_shiftReg_40_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(141.235 11.49 141.365 11.64)
MU9413/5/reg_r_shiftReg_40_/8 G_DG U9413/5/265 U9413/5/reg_r_shiftReg_40_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(141.715 11.49 141.845 11.64)
MU9413/5/reg_r_shiftReg_40_/9 U9413/5/reg_r_shiftReg_40_/9 U9413/5/268 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(142.805 11.49 142.935 11.64)
MU9413/5/reg_r_shiftReg_40_/10 U9413/5/reg_r_shiftReg_40_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_40_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(143.315 11.49 143.445 11.64)
MU9413/5/reg_r_shiftReg_40_/11 U9413/5/271 U9413/5/265 U9413/5/reg_r_shiftReg_40_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(143.735 11.49 143.865 11.64)
MU9413/5/reg_r_shiftReg_40_/12 U9413/5/272 U9413/5/271 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(144.825 11.49 144.955 11.64)
MU9413/5/reg_r_shiftReg_40_/13 U9413/5/273 U9413/5/264 U9413/5/271 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(146.185 11.49 146.315 11.64)
MU9413/5/reg_r_shiftReg_40_/14 U9413/5/reg_r_shiftReg_40_/14 U9413/5/CLB U9413/5/273 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(146.765 11.49 146.895 11.64)
MU9413/5/reg_r_shiftReg_40_/15 G_DG U9413/5/272 U9413/5/reg_r_shiftReg_40_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(147.075 11.49 147.205 11.64)
MU9413/5/reg_r_shiftReg_40_/16 addr[7] U9413/5/273 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(148.165 11.49 148.295 11.64)
MU9413/5/reg_r_shiftReg_40_/17 U9413/5/reg_r_shiftReg_40_/QB U9413/5/272 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(149.255 11.49 149.385 11.64)
MU9413/5/ix1776/1 G_DG U9413/SEL U9413/5/260 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(132.03 11.49 132.16 11.64)
MU9413/5/ix1776/2 U9413/5/ix1776/3 U9413/5/260 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(132.61 11.49 132.74 11.64)
MU9413/5/ix1776/3 U9413/5/262 addr[7] U9413/5/ix1776/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(133.19 11.49 133.32 11.64)
MU9413/5/ix1776/4 U9413/5/ix1776/5 addr[6] U9413/5/262 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(133.77 11.49 133.9 11.64)
MU9413/5/ix1776/5 G_DG U9413/SEL U9413/5/ix1776/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(134.35 11.49 134.48 11.64)
MU9413/5/ix1776/6 U9413/5/DATA U9413/5/262 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(134.93 11.49 135.06 11.64)
MU9413/5/ix1766/1 G_DG U9413/6/SEL U9413/5/253 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(127.95 11.49 128.08 11.64)
MU9413/5/ix1766/2 U9413/5/ix1766/3 U9413/5/253 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(128.53 11.49 128.66 11.64)
MU9413/5/ix1766/3 U9413/5/255 addr[6] U9413/5/ix1766/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(129.11 11.49 129.24 11.64)
MU9413/5/ix1766/4 U9413/5/ix1766/5 addr[5] U9413/5/255 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(129.69 11.49 129.82 11.64)
MU9413/5/ix1766/5 G_DG U9413/6/SEL U9413/5/ix1766/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(130.27 11.49 130.4 11.64)
MU9413/5/ix1766/6 U9413/5/ix1766/OUT U9413/5/255 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(130.85 11.49 130.98 11.64)
MU9413/5/reg_r_shiftReg_39_/1 G_DG U9413/5/CLK U9413/5/239 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(113.625 11.49 113.755 11.64)
MU9413/5/reg_r_shiftReg_39_/2 U9413/5/240 U9413/5/239 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(114.205 11.49 114.335 11.64)
MU9413/5/reg_r_shiftReg_39_/3 U9413/5/reg_r_shiftReg_39_/4 U9413/5/ix1766/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(115.295 11.49 115.425 11.64)
MU9413/5/reg_r_shiftReg_39_/4 U9413/5/243 U9413/5/239 U9413/5/reg_r_shiftReg_39_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(115.81 11.49 115.94 11.64)
MU9413/5/reg_r_shiftReg_39_/5 U9413/5/244 U9413/5/243 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(116.9 11.49 117.03 11.64)
MU9413/5/reg_r_shiftReg_39_/6 U9413/5/reg_r_shiftReg_39_/7 U9413/5/CLB U9413/5/243 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(118.27 11.49 118.4 11.64)
MU9413/5/reg_r_shiftReg_39_/7 U9413/5/reg_r_shiftReg_39_/8 U9413/5/244 U9413/5/reg_r_shiftReg_39_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(118.75 11.49 118.88 11.64)
MU9413/5/reg_r_shiftReg_39_/8 G_DG U9413/5/240 U9413/5/reg_r_shiftReg_39_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(119.23 11.49 119.36 11.64)
MU9413/5/reg_r_shiftReg_39_/9 U9413/5/reg_r_shiftReg_39_/9 U9413/5/244 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(120.32 11.49 120.45 11.64)
MU9413/5/reg_r_shiftReg_39_/10 U9413/5/reg_r_shiftReg_39_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_39_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(120.83 11.49 120.96 11.64)
MU9413/5/reg_r_shiftReg_39_/11 U9413/5/247 U9413/5/240 U9413/5/reg_r_shiftReg_39_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(121.25 11.49 121.38 11.64)
MU9413/5/reg_r_shiftReg_39_/12 U9413/5/248 U9413/5/247 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(122.34 11.49 122.47 11.64)
MU9413/5/reg_r_shiftReg_39_/13 U9413/5/249 U9413/5/239 U9413/5/247 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(123.7 11.49 123.83 11.64)
MU9413/5/reg_r_shiftReg_39_/14 U9413/5/reg_r_shiftReg_39_/14 U9413/5/CLB U9413/5/249 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(124.28 11.49 124.41 11.64)
MU9413/5/reg_r_shiftReg_39_/15 G_DG U9413/5/248 U9413/5/reg_r_shiftReg_39_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(124.59 11.49 124.72 11.64)
MU9413/5/reg_r_shiftReg_39_/16 addr[6] U9413/5/249 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(125.68 11.49 125.81 11.64)
MU9413/5/reg_r_shiftReg_39_/17 U9413/5/reg_r_shiftReg_39_/QB U9413/5/248 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(126.77 11.49 126.9 11.64)
MU9413/5/reg_r_shiftReg_3_/1 G_DG U9413/5/CLK U9413/5/226 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(99.3 11.49 99.43 11.64)
MU9413/5/reg_r_shiftReg_3_/2 U9413/5/227 U9413/5/226 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(99.88 11.49 100.01 11.64)
MU9413/5/reg_r_shiftReg_3_/3 U9413/5/reg_r_shiftReg_3_/4 U9413/ix1786\Cross G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(100.97 11.49 101.1 11.64)
MU9413/5/reg_r_shiftReg_3_/4 U9413/5/230 U9413/5/226 U9413/5/reg_r_shiftReg_3_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(101.485 11.49 101.615 11.64)
MU9413/5/reg_r_shiftReg_3_/5 U9413/5/231 U9413/5/230 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(102.575 11.49 102.705 11.64)
MU9413/5/reg_r_shiftReg_3_/6 U9413/5/reg_r_shiftReg_3_/7 U9413/5/CLB U9413/5/230 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(103.945 11.49 104.075 11.64)
MU9413/5/reg_r_shiftReg_3_/7 U9413/5/reg_r_shiftReg_3_/8 U9413/5/231 U9413/5/reg_r_shiftReg_3_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(104.425 11.49 104.555 11.64)
MU9413/5/reg_r_shiftReg_3_/8 G_DG U9413/5/227 U9413/5/reg_r_shiftReg_3_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(104.905 11.49 105.035 11.64)
MU9413/5/reg_r_shiftReg_3_/9 U9413/5/reg_r_shiftReg_3_/9 U9413/5/231 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(105.995 11.49 106.125 11.64)
MU9413/5/reg_r_shiftReg_3_/10 U9413/5/reg_r_shiftReg_3_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_3_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(106.505 11.49 106.635 11.64)
MU9413/5/reg_r_shiftReg_3_/11 U9413/5/234 U9413/5/227 U9413/5/reg_r_shiftReg_3_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(106.925 11.49 107.055 11.64)
MU9413/5/reg_r_shiftReg_3_/12 U9413/5/235 U9413/5/234 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(108.015 11.49 108.145 11.64)
MU9413/5/reg_r_shiftReg_3_/13 U9413/5/236 U9413/5/226 U9413/5/234 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(109.375 11.49 109.505 11.64)
MU9413/5/reg_r_shiftReg_3_/14 U9413/5/reg_r_shiftReg_3_/14 U9413/5/CLB U9413/5/236 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(109.955 11.49 110.085 11.64)
MU9413/5/reg_r_shiftReg_3_/15 G_DG U9413/5/235 U9413/5/reg_r_shiftReg_3_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(110.265 11.49 110.395 11.64)
MU9413/5/reg_r_shiftReg_3_/16 wrData[2] U9413/5/236 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(111.355 11.49 111.485 11.64)
MU9413/5/reg_r_shiftReg_3_/17 U9413/5/reg_r_shiftReg_3_/QB U9413/5/235 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(112.445 11.49 112.575 11.64)
MU9413/5/ix47/1 U9413/D ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(97.54 11.49 97.67 11.64)
MU9413/5/ix47/2 G_DG U9413/6/SEL U9413/D G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(98.12 11.49 98.25 11.64)
MU9413/5/reg_r_shiftReg_35_/1 G_DG U9413/5/CLK U9413/5/209 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(83.215 11.49 83.345 11.64)
MU9413/5/reg_r_shiftReg_35_/2 U9413/5/210 U9413/5/209 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(83.795 11.49 83.925 11.64)
MU9413/5/reg_r_shiftReg_35_/3 U9413/5/reg_r_shiftReg_35_/4 U9413/5/reg_r_shiftReg_35_/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(84.885 11.49 85.015 11.64)
MU9413/5/reg_r_shiftReg_35_/4 U9413/5/213 U9413/5/209 U9413/5/reg_r_shiftReg_35_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(85.4 11.49 85.53 11.64)
MU9413/5/reg_r_shiftReg_35_/5 U9413/5/214 U9413/5/213 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(86.49 11.49 86.62 11.64)
MU9413/5/reg_r_shiftReg_35_/6 U9413/5/reg_r_shiftReg_35_/7 U9413/5/CLB U9413/5/213 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(87.86 11.49 87.99 11.64)
MU9413/5/reg_r_shiftReg_35_/7 U9413/5/reg_r_shiftReg_35_/8 U9413/5/214 U9413/5/reg_r_shiftReg_35_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(88.34 11.49 88.47 11.64)
MU9413/5/reg_r_shiftReg_35_/8 G_DG U9413/5/210 U9413/5/reg_r_shiftReg_35_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(88.82 11.49 88.95 11.64)
MU9413/5/reg_r_shiftReg_35_/9 U9413/5/reg_r_shiftReg_35_/9 U9413/5/214 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(89.91 11.49 90.04 11.64)
MU9413/5/reg_r_shiftReg_35_/10 U9413/5/reg_r_shiftReg_35_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_35_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(90.42 11.49 90.55 11.64)
MU9413/5/reg_r_shiftReg_35_/11 U9413/5/217 U9413/5/210 U9413/5/reg_r_shiftReg_35_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(90.84 11.49 90.97 11.64)
MU9413/5/reg_r_shiftReg_35_/12 U9413/5/218 U9413/5/217 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(91.93 11.49 92.06 11.64)
MU9413/5/reg_r_shiftReg_35_/13 U9413/5/219 U9413/5/209 U9413/5/217 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(93.29 11.49 93.42 11.64)
MU9413/5/reg_r_shiftReg_35_/14 U9413/5/reg_r_shiftReg_35_/14 U9413/5/CLB U9413/5/219 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(93.87 11.49 94 11.64)
MU9413/5/reg_r_shiftReg_35_/15 G_DG U9413/5/218 U9413/5/reg_r_shiftReg_35_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(94.18 11.49 94.31 11.64)
MU9413/5/reg_r_shiftReg_35_/16 addr[2] U9413/5/219 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(95.27 11.49 95.4 11.64)
MU9413/5/reg_r_shiftReg_35_/17 U9413/5/reg_r_shiftReg_35_/QB U9413/5/218 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(96.36 11.49 96.49 11.64)
MU9413/5/reg_r_shiftReg_8_/1 G_DG U9413/5/CLK U9413/5/196 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(68.89 11.49 69.02 11.64)
MU9413/5/reg_r_shiftReg_8_/2 U9413/5/197 U9413/5/196 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(69.47 11.49 69.6 11.64)
MU9413/5/reg_r_shiftReg_8_/3 U9413/5/reg_r_shiftReg_8_/4 U9413/4/ix145/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(70.56 11.49 70.69 11.64)
MU9413/5/reg_r_shiftReg_8_/4 U9413/5/200 U9413/5/196 U9413/5/reg_r_shiftReg_8_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(71.075 11.49 71.205 11.64)
MU9413/5/reg_r_shiftReg_8_/5 U9413/5/201 U9413/5/200 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(72.165 11.49 72.295 11.64)
MU9413/5/reg_r_shiftReg_8_/6 U9413/5/reg_r_shiftReg_8_/7 U9413/5/CLB U9413/5/200 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(73.535 11.49 73.665 11.64)
MU9413/5/reg_r_shiftReg_8_/7 U9413/5/reg_r_shiftReg_8_/8 U9413/5/201 U9413/5/reg_r_shiftReg_8_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(74.015 11.49 74.145 11.64)
MU9413/5/reg_r_shiftReg_8_/8 G_DG U9413/5/197 U9413/5/reg_r_shiftReg_8_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(74.495 11.49 74.625 11.64)
MU9413/5/reg_r_shiftReg_8_/9 U9413/5/reg_r_shiftReg_8_/9 U9413/5/201 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(75.585 11.49 75.715 11.64)
MU9413/5/reg_r_shiftReg_8_/10 U9413/5/reg_r_shiftReg_8_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_8_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(76.095 11.49 76.225 11.64)
MU9413/5/reg_r_shiftReg_8_/11 U9413/5/204 U9413/5/197 U9413/5/reg_r_shiftReg_8_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(76.515 11.49 76.645 11.64)
MU9413/5/reg_r_shiftReg_8_/12 U9413/5/205 U9413/5/204 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(77.605 11.49 77.735 11.64)
MU9413/5/reg_r_shiftReg_8_/13 U9413/5/206 U9413/5/196 U9413/5/204 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(78.965 11.49 79.095 11.64)
MU9413/5/reg_r_shiftReg_8_/14 U9413/5/reg_r_shiftReg_8_/14 U9413/5/CLB U9413/5/206 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(79.545 11.49 79.675 11.64)
MU9413/5/reg_r_shiftReg_8_/15 G_DG U9413/5/205 U9413/5/reg_r_shiftReg_8_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(79.855 11.49 79.985 11.64)
MU9413/5/reg_r_shiftReg_8_/16 wrData[7] U9413/5/206 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(80.945 11.49 81.075 11.64)
MU9413/5/reg_r_shiftReg_8_/17 U9413/5/reg_r_shiftReg_8_/QB U9413/5/205 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(82.035 11.49 82.165 11.64)
MU9413/5/reg_r_shiftReg_13_/1 G_DG U9413/5/CLK U9413/5/183 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(54.565 11.49 54.695 11.64)
MU9413/5/reg_r_shiftReg_13_/2 U9413/5/184 U9413/5/183 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(55.145 11.49 55.275 11.64)
MU9413/5/reg_r_shiftReg_13_/3 U9413/5/reg_r_shiftReg_13_/4 U9413/4/ix205/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(56.235 11.49 56.365 11.64)
MU9413/5/reg_r_shiftReg_13_/4 U9413/5/187 U9413/5/183 U9413/5/reg_r_shiftReg_13_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(56.75 11.49 56.88 11.64)
MU9413/5/reg_r_shiftReg_13_/5 U9413/5/188 U9413/5/187 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(57.84 11.49 57.97 11.64)
MU9413/5/reg_r_shiftReg_13_/6 U9413/5/reg_r_shiftReg_13_/7 U9413/5/CLB U9413/5/187 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(59.21 11.49 59.34 11.64)
MU9413/5/reg_r_shiftReg_13_/7 U9413/5/reg_r_shiftReg_13_/8 U9413/5/188 U9413/5/reg_r_shiftReg_13_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(59.69 11.49 59.82 11.64)
MU9413/5/reg_r_shiftReg_13_/8 G_DG U9413/5/184 U9413/5/reg_r_shiftReg_13_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(60.17 11.49 60.3 11.64)
MU9413/5/reg_r_shiftReg_13_/9 U9413/5/reg_r_shiftReg_13_/9 U9413/5/188 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(61.26 11.49 61.39 11.64)
MU9413/5/reg_r_shiftReg_13_/10 U9413/5/reg_r_shiftReg_13_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_13_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(61.77 11.49 61.9 11.64)
MU9413/5/reg_r_shiftReg_13_/11 U9413/5/191 U9413/5/184 U9413/5/reg_r_shiftReg_13_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(62.19 11.49 62.32 11.64)
MU9413/5/reg_r_shiftReg_13_/12 U9413/5/192 U9413/5/191 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(63.28 11.49 63.41 11.64)
MU9413/5/reg_r_shiftReg_13_/13 U9413/5/193 U9413/5/183 U9413/5/191 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(64.64 11.49 64.77 11.64)
MU9413/5/reg_r_shiftReg_13_/14 U9413/5/reg_r_shiftReg_13_/14 U9413/5/CLB U9413/5/193 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(65.22 11.49 65.35 11.64)
MU9413/5/reg_r_shiftReg_13_/15 G_DG U9413/5/192 U9413/5/reg_r_shiftReg_13_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(65.53 11.49 65.66 11.64)
MU9413/5/reg_r_shiftReg_13_/16 wrData[12] U9413/5/193 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(66.62 11.49 66.75 11.64)
MU9413/5/reg_r_shiftReg_13_/17 U9413/5/reg_r_shiftReg_13_/QB U9413/5/192 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(67.71 11.49 67.84 11.64)
MU9413/5/ix1826/1 G_DG U9413/SEL U9413/5/176 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(50.485 11.49 50.615 11.64)
MU9413/5/ix1826/2 U9413/5/ix1826/3 U9413/5/176 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(51.065 11.49 51.195 11.64)
MU9413/5/ix1826/3 U9413/5/178 cmd[0] U9413/5/ix1826/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(51.645 11.49 51.775 11.64)
MU9413/5/ix1826/4 U9413/5/ix1826/5 addr[11] U9413/5/178 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(52.225 11.49 52.355 11.64)
MU9413/5/ix1826/5 G_DG U9413/SEL U9413/5/ix1826/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(52.805 11.49 52.935 11.64)
MU9413/5/ix1826/6 U9413/5/ix1826/OUT U9413/5/178 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(53.385 11.49 53.515 11.64)
MU9413/5/reg_r_shiftReg_15_/1 G_DG U9413/5/CLK U9413/5/162 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(36.16 11.49 36.29 11.64)
MU9413/5/reg_r_shiftReg_15_/2 U9413/5/163 U9413/5/162 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(36.74 11.49 36.87 11.64)
MU9413/5/reg_r_shiftReg_15_/3 U9413/5/reg_r_shiftReg_15_/4 U9413/4/ix229/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(37.83 11.49 37.96 11.64)
MU9413/5/reg_r_shiftReg_15_/4 U9413/5/166 U9413/5/162 U9413/5/reg_r_shiftReg_15_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(38.345 11.49 38.475 11.64)
MU9413/5/reg_r_shiftReg_15_/5 U9413/5/167 U9413/5/166 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(39.435 11.49 39.565 11.64)
MU9413/5/reg_r_shiftReg_15_/6 U9413/5/reg_r_shiftReg_15_/7 U9413/5/CLB U9413/5/166 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(40.805 11.49 40.935 11.64)
MU9413/5/reg_r_shiftReg_15_/7 U9413/5/reg_r_shiftReg_15_/8 U9413/5/167 U9413/5/reg_r_shiftReg_15_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(41.285 11.49 41.415 11.64)
MU9413/5/reg_r_shiftReg_15_/8 G_DG U9413/5/163 U9413/5/reg_r_shiftReg_15_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(41.765 11.49 41.895 11.64)
MU9413/5/reg_r_shiftReg_15_/9 U9413/5/reg_r_shiftReg_15_/9 U9413/5/167 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(42.855 11.49 42.985 11.64)
MU9413/5/reg_r_shiftReg_15_/10 U9413/5/reg_r_shiftReg_15_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_15_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(43.365 11.49 43.495 11.64)
MU9413/5/reg_r_shiftReg_15_/11 U9413/5/170 U9413/5/163 U9413/5/reg_r_shiftReg_15_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(43.785 11.49 43.915 11.64)
MU9413/5/reg_r_shiftReg_15_/12 U9413/5/171 U9413/5/170 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(44.875 11.49 45.005 11.64)
MU9413/5/reg_r_shiftReg_15_/13 U9413/5/172 U9413/5/162 U9413/5/170 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(46.235 11.49 46.365 11.64)
MU9413/5/reg_r_shiftReg_15_/14 U9413/5/reg_r_shiftReg_15_/14 U9413/5/CLB U9413/5/172 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(46.815 11.49 46.945 11.64)
MU9413/5/reg_r_shiftReg_15_/15 G_DG U9413/5/171 U9413/5/reg_r_shiftReg_15_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(47.125 11.49 47.255 11.64)
MU9413/5/reg_r_shiftReg_15_/16 wrData[14] U9413/5/172 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(48.215 11.49 48.345 11.64)
MU9413/5/reg_r_shiftReg_15_/17 U9413/5/reg_r_shiftReg_15_/QB U9413/5/171 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(49.305 11.49 49.435 11.64)
MU9413/5/reg_r_shiftReg_0_/1 G_DG U9413/5/CLK U9413/5/149 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(21.835 11.49 21.965 11.64)
MU9413/5/reg_r_shiftReg_0_/2 U9413/5/150 U9413/5/149 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(22.415 11.49 22.545 11.64)
MU9413/5/reg_r_shiftReg_0_/3 U9413/5/reg_r_shiftReg_0_/4 U9413/5/reg_r_shiftReg_0_/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(23.505 11.49 23.635 11.64)
MU9413/5/reg_r_shiftReg_0_/4 U9413/5/153 U9413/5/149 U9413/5/reg_r_shiftReg_0_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(24.02 11.49 24.15 11.64)
MU9413/5/reg_r_shiftReg_0_/5 U9413/5/154 U9413/5/153 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(25.11 11.49 25.24 11.64)
MU9413/5/reg_r_shiftReg_0_/6 U9413/5/reg_r_shiftReg_0_/7 U9413/5/CLB U9413/5/153 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(26.48 11.49 26.61 11.64)
MU9413/5/reg_r_shiftReg_0_/7 U9413/5/reg_r_shiftReg_0_/8 U9413/5/154 U9413/5/reg_r_shiftReg_0_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(26.96 11.49 27.09 11.64)
MU9413/5/reg_r_shiftReg_0_/8 G_DG U9413/5/150 U9413/5/reg_r_shiftReg_0_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(27.44 11.49 27.57 11.64)
MU9413/5/reg_r_shiftReg_0_/9 U9413/5/reg_r_shiftReg_0_/9 U9413/5/154 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(28.53 11.49 28.66 11.64)
MU9413/5/reg_r_shiftReg_0_/10 U9413/5/reg_r_shiftReg_0_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_0_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(29.04 11.49 29.17 11.64)
MU9413/5/reg_r_shiftReg_0_/11 U9413/5/157 U9413/5/150 U9413/5/reg_r_shiftReg_0_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(29.46 11.49 29.59 11.64)
MU9413/5/reg_r_shiftReg_0_/12 U9413/5/158 U9413/5/157 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(30.55 11.49 30.68 11.64)
MU9413/5/reg_r_shiftReg_0_/13 U9413/5/159 U9413/5/149 U9413/5/157 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(31.91 11.49 32.04 11.64)
MU9413/5/reg_r_shiftReg_0_/14 U9413/5/reg_r_shiftReg_0_/14 U9413/5/CLB U9413/5/159 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(32.49 11.49 32.62 11.64)
MU9413/5/reg_r_shiftReg_0_/15 G_DG U9413/5/158 U9413/5/reg_r_shiftReg_0_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(32.8 11.49 32.93 11.64)
MU9413/5/reg_r_shiftReg_0_/16 U9413/4/ix2251/A U9413/5/159 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(33.89 11.49 34.02 11.64)
MU9413/5/reg_r_shiftReg_0_/17 U9413/5/reg_r_shiftReg_0_/QB U9413/5/158 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(34.98 11.49 35.11 11.64)
MU9413/5/ix2272/1 G_DG U9413/5/ix2272/A U9413/5/147 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(20.075 11.49 20.205 11.64)
MU9413/5/ix2272/2 U9413/SEL U9413/5/147 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(20.655 11.49 20.785 11.64)
MU9413/5/ix2298/1 G_DG U9413/5/ix2272/A U9413/5/144 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(18.315 11.49 18.445 11.64)
MU9413/5/ix2298/2 U9413/6/SEL U9413/5/144 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(18.895 11.49 19.025 11.64)
MU9413/5/reg_r_state/1 G_DG U9413/5/CLK U9413/5/131 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(3.99 11.49 4.12 11.64)
MU9413/5/reg_r_state/2 U9413/5/132 U9413/5/131 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(4.57 11.49 4.7 11.64)
MU9413/5/reg_r_state/3 U9413/5/reg_r_state/4 U9413/5/ix25/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(5.66 11.49 5.79 11.64)
MU9413/5/reg_r_state/4 U9413/5/135 U9413/5/131 U9413/5/reg_r_state/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(6.175 11.49 6.305 11.64)
MU9413/5/reg_r_state/5 U9413/5/136 U9413/5/135 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(7.265 11.49 7.395 11.64)
MU9413/5/reg_r_state/6 U9413/5/reg_r_state/7 U9413/5/CLB U9413/5/135 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(8.635 11.49 8.765 11.64)
MU9413/5/reg_r_state/7 U9413/5/reg_r_state/8 U9413/5/136 U9413/5/reg_r_state/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(9.115 11.49 9.245 11.64)
MU9413/5/reg_r_state/8 G_DG U9413/5/132 U9413/5/reg_r_state/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(9.595 11.49 9.725 11.64)
MU9413/5/reg_r_state/9 U9413/5/reg_r_state/9 U9413/5/136 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(10.685 11.49 10.815 11.64)
MU9413/5/reg_r_state/10 U9413/5/reg_r_state/10 U9413/5/CLB U9413/5/reg_r_state/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(11.195 11.49 11.325 11.64)
MU9413/5/reg_r_state/11 U9413/5/139 U9413/5/132 U9413/5/reg_r_state/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(11.615 11.49 11.745 11.64)
MU9413/5/reg_r_state/12 U9413/5/140 U9413/5/139 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(12.705 11.49 12.835 11.64)
MU9413/5/reg_r_state/13 U9413/5/141 U9413/5/131 U9413/5/139 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(14.065 11.49 14.195 11.64)
MU9413/5/reg_r_state/14 U9413/5/reg_r_state/14 U9413/5/CLB U9413/5/141 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(14.645 11.49 14.775 11.64)
MU9413/5/reg_r_state/15 G_DG U9413/5/140 U9413/5/reg_r_state/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(14.955 11.49 15.085 11.64)
MU9413/5/reg_r_state/16 U9413/5/ix39/B U9413/5/141 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(16.045 11.49 16.175 11.64)
MU9413/5/reg_r_state/17 U9413/QB U9413/5/140 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(17.135 11.49 17.265 11.64)
MU9413/5/ix39/1 U9413/5/ix39/1 U9413/5/ix2198/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(2.23 11.49 2.36 11.64)
MU9413/5/ix39/2 U9413/4/ix2276/A U9413/5/ix39/B U9413/5/ix39/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(2.81 11.49 2.94 11.64)
MU9413/5/ix9_0_XREP9/1 U9413/5/ix9_0_XREP9/1 exec G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(0.47 11.49 0.6 11.64)
MU9413/5/ix9_0_XREP9/2 U9413/5/ix2272/A U9413/5/C U9413/5/ix9_0_XREP9/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(1.05 11.49 1.18 11.64)
MU9413/5/ix2198/1 U9413/5/ix2198/1 U9413/6/QB G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-1.88 11.49 -1.75 11.64)
MU9413/5/ix2198/2 U9413/5/ix2198/3 U9413/5/ix2004/OUT U9413/5/ix2198/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=3.45e-014 pd=6.1e-007 ps=6e-007 nrd=1.53333 nrs=1.5  $(-1.3 11.49 -1.17 11.64)
MU9413/5/ix2198/3 U9413/5/ix2198/OUT U9413/5/C U9413/5/ix2198/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.45e-014 ad=1.3425e-013 pd=1.57e-006 ps=6.1e-007 nrd=5.96667 nrs=1.53333  $(-0.71 11.49 -0.58 11.64)
MU9413/5/ix2198/4 U9413/5/ix2198/OUT U9413/6/QB G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=1.365e-013 ad=7.8e-014 pd=8.4e-007 ps=1.53e-006 nrd=1.15385 nrs=2.01923  $(-1.88 13.22 -1.75 13.48)
MU9413/5/ix2198/5 G_DS U9413/5/ix2004/OUT U9413/5/ix2198/OUT G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.8e-014 ad=7.93e-014 pd=8.5e-007 ps=8.4e-007 nrd=1.17308 nrs=1.15385  $(-1.3 13.22 -1.17 13.48)
MU9413/5/ix2198/6 U9413/5/ix2198/OUT U9413/5/C G_DS G_DS pch sa=-1 sb=-1 w=2.6e-007 l=1.3e-007 as=7.93e-014 ad=1.365e-013 pd=1.53e-006 ps=8.5e-007 nrd=2.01923 nrs=1.17308  $(-0.71 13.22 -0.58 13.48)
MU9413/5/ix25/1 G_DG U9413/QB U9413/5/118 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-5.96 11.49 -5.83 11.64)
MU9413/5/ix25/2 U9413/5/ix25/3 U9413/5/118 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-5.38 11.49 -5.25 11.64)
MU9413/5/ix25/3 U9413/5/120 U9413/5/ix2004/OUT U9413/5/ix25/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-4.8 11.49 -4.67 11.64)
MU9413/5/ix25/4 U9413/5/ix25/5 U9413/4/ix2251/A U9413/5/120 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-4.22 11.49 -4.09 11.64)
MU9413/5/ix25/5 G_DG U9413/QB U9413/5/ix25/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-3.64 11.49 -3.51 11.64)
MU9413/5/ix25/6 U9413/5/ix25/OUT U9413/5/120 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-3.06 11.49 -2.93 11.64)
MU9413/5/ix2004/1 U9413/5/ix2004/OUT ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-7.14 11.49 -7.01 11.64)
MU9413/5/ix55/1 U9413/3/ix2292/A U9413/5/ix1896/B G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-9.48 11.49 -9.35 11.64)
MU9413/5/ix55/2 G_DG U9413/5/ix2004/OUT U9413/3/ix2292/A G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=7.275e-014 pd=8.6e-007 ps=8.6e-007 nrd=3.23333 nrs=3.23333  $(-8.9 11.49 -8.77 11.64)
MU9413/5/ix55/3 U9413/3/ix2292/A U9413/5/ix489/B G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-8.32 11.49 -8.19 11.64)
MU9413/5/reg_r_state_0_XREP7/1 G_DG U9413/5/CLK U9413/5/96 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-23.805 11.49 -23.675 11.64)
MU9413/5/reg_r_state_0_XREP7/2 U9413/5/97 U9413/5/96 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-23.225 11.49 -23.095 11.64)
MU9413/5/reg_r_state_0_XREP7/3 U9413/5/reg_r_state_0_XREP7/4 U9413/5/ix25/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-22.135 11.49 -22.005 11.64)
MU9413/5/reg_r_state_0_XREP7/4 U9413/5/100 U9413/5/96 U9413/5/reg_r_state_0_XREP7/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-21.62 11.49 -21.49 11.64)
MU9413/5/reg_r_state_0_XREP7/5 U9413/5/101 U9413/5/100 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-20.53 11.49 -20.4 11.64)
MU9413/5/reg_r_state_0_XREP7/6 U9413/5/reg_r_state_0_XREP7/7 U9413/5/CLB U9413/5/100 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-19.16 11.49 -19.03 11.64)
MU9413/5/reg_r_state_0_XREP7/7 U9413/5/reg_r_state_0_XREP7/8 U9413/5/101 U9413/5/reg_r_state_0_XREP7/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-18.68 11.49 -18.55 11.64)
MU9413/5/reg_r_state_0_XREP7/8 G_DG U9413/5/97 U9413/5/reg_r_state_0_XREP7/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-18.2 11.49 -18.07 11.64)
MU9413/5/reg_r_state_0_XREP7/9 U9413/5/reg_r_state_0_XREP7/9 U9413/5/101 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-17.11 11.49 -16.98 11.64)
MU9413/5/reg_r_state_0_XREP7/10 U9413/5/reg_r_state_0_XREP7/10 U9413/5/CLB U9413/5/reg_r_state_0_XREP7/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-16.6 11.49 -16.47 11.64)
MU9413/5/reg_r_state_0_XREP7/11 U9413/5/104 U9413/5/97 U9413/5/reg_r_state_0_XREP7/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-16.18 11.49 -16.05 11.64)
MU9413/5/reg_r_state_0_XREP7/12 U9413/5/105 U9413/5/104 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-15.09 11.49 -14.96 11.64)
MU9413/5/reg_r_state_0_XREP7/13 U9413/5/106 U9413/5/96 U9413/5/104 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-13.73 11.49 -13.6 11.64)
MU9413/5/reg_r_state_0_XREP7/14 U9413/5/reg_r_state_0_XREP7/14 U9413/5/CLB U9413/5/106 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-13.15 11.49 -13.02 11.64)
MU9413/5/reg_r_state_0_XREP7/15 G_DG U9413/5/105 U9413/5/reg_r_state_0_XREP7/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-12.84 11.49 -12.71 11.64)
MU9413/5/reg_r_state_0_XREP7/16 U9413/5/C U9413/5/106 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-11.75 11.49 -11.62 11.64)
MU9413/5/reg_r_state_0_XREP7/17 U9413/5/ix489/B U9413/5/105 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-10.66 11.49 -10.53 11.64)
MU9413/5/ix9/1 U9413/5/ix9/1 exec G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=3.375e-014 pd=6e-007 ps=1.57e-006 nrd=1.5 nrs=5.96667  $(-25.565 11.49 -25.435 11.64)
MU9413/5/ix9/2 U9413/4/ix2270/A U9413/5/C U9413/5/ix9/1 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=1.3425e-013 pd=1.57e-006 ps=6e-007 nrd=5.96667 nrs=1.5  $(-24.985 11.49 -24.855 11.64)
MU9413/5/ix2274/1 G_DG U9413/4/ix2270/A U9413/5/91 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-27.325 11.49 -27.195 11.64)
MU9413/5/ix2274/2 U9413/5/ix1876/SEL U9413/5/91 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-26.745 11.49 -26.615 11.64)
MU9413/5/reg_r_shiftReg_52_/1 G_DG U9413/5/CLK U9413/5/77 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-41.65 11.49 -41.52 11.64)
MU9413/5/reg_r_shiftReg_52_/2 U9413/5/78 U9413/5/77 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-41.07 11.49 -40.94 11.64)
MU9413/5/reg_r_shiftReg_52_/3 U9413/5/reg_r_shiftReg_52_/4 U9413/5/ix1896/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-39.98 11.49 -39.85 11.64)
MU9413/5/reg_r_shiftReg_52_/4 U9413/5/81 U9413/5/77 U9413/5/reg_r_shiftReg_52_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-39.465 11.49 -39.335 11.64)
MU9413/5/reg_r_shiftReg_52_/5 U9413/5/82 U9413/5/81 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-38.375 11.49 -38.245 11.64)
MU9413/5/reg_r_shiftReg_52_/6 U9413/5/reg_r_shiftReg_52_/7 U9413/5/CLB U9413/5/81 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-37.005 11.49 -36.875 11.64)
MU9413/5/reg_r_shiftReg_52_/7 U9413/5/reg_r_shiftReg_52_/8 U9413/5/82 U9413/5/reg_r_shiftReg_52_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-36.525 11.49 -36.395 11.64)
MU9413/5/reg_r_shiftReg_52_/8 G_DG U9413/5/78 U9413/5/reg_r_shiftReg_52_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-36.045 11.49 -35.915 11.64)
MU9413/5/reg_r_shiftReg_52_/9 U9413/5/reg_r_shiftReg_52_/9 U9413/5/82 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-34.955 11.49 -34.825 11.64)
MU9413/5/reg_r_shiftReg_52_/10 U9413/5/reg_r_shiftReg_52_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_52_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-34.445 11.49 -34.315 11.64)
MU9413/5/reg_r_shiftReg_52_/11 U9413/5/85 U9413/5/78 U9413/5/reg_r_shiftReg_52_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-34.025 11.49 -33.895 11.64)
MU9413/5/reg_r_shiftReg_52_/12 U9413/5/86 U9413/5/85 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-32.935 11.49 -32.805 11.64)
MU9413/5/reg_r_shiftReg_52_/13 U9413/5/87 U9413/5/77 U9413/5/85 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-31.575 11.49 -31.445 11.64)
MU9413/5/reg_r_shiftReg_52_/14 U9413/5/reg_r_shiftReg_52_/14 U9413/5/CLB U9413/5/87 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-30.995 11.49 -30.865 11.64)
MU9413/5/reg_r_shiftReg_52_/15 G_DG U9413/5/86 U9413/5/reg_r_shiftReg_52_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-30.685 11.49 -30.555 11.64)
MU9413/5/reg_r_shiftReg_52_/16 U9413/5/ix1896/B U9413/5/87 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-29.595 11.49 -29.465 11.64)
MU9413/5/reg_r_shiftReg_52_/17 U9413/5/ix489/C U9413/5/86 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-28.505 11.49 -28.375 11.64)
MU9413/5/ix489/1 U9413/5/ix1916/SEL exec G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-43.99 11.49 -43.86 11.64)
MU9413/5/ix489/2 G_DG U9413/5/ix489/B U9413/5/ix1916/SEL G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=7.275e-014 pd=8.6e-007 ps=8.6e-007 nrd=3.23333 nrs=3.23333  $(-43.41 11.49 -43.28 11.64)
MU9413/5/ix489/3 U9413/5/ix1916/SEL U9413/5/ix489/C G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-42.83 11.49 -42.7 11.64)
MU9413/5/ix1896/1 G_DG U9413/5/ix1876/SEL U9413/5/64 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-48.07 11.49 -47.94 11.64)
MU9413/5/ix1896/2 U9413/5/ix1896/3 U9413/5/64 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-47.49 11.49 -47.36 11.64)
MU9413/5/ix1896/3 U9413/5/66 U9413/5/ix1896/B U9413/5/ix1896/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-46.91 11.49 -46.78 11.64)
MU9413/5/ix1896/4 U9413/5/ix1896/5 cmd[6] U9413/5/66 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-46.33 11.49 -46.2 11.64)
MU9413/5/ix1896/5 G_DG U9413/5/ix1876/SEL U9413/5/ix1896/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-45.75 11.49 -45.62 11.64)
MU9413/5/ix1896/6 U9413/5/ix1896/OUT U9413/5/66 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-45.17 11.49 -45.04 11.64)
MU9413/5/ix1916/1 G_DG U9413/5/ix1916/SEL U9413/5/56 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-52.15 11.49 -52.02 11.64)
MU9413/5/ix1916/2 U9413/5/ix1916/3 U9413/5/56 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-51.57 11.49 -51.44 11.64)
MU9413/5/ix1916/3 U9413/5/58 readL U9413/5/ix1916/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-50.99 11.49 -50.86 11.64)
MU9413/5/ix1916/4 U9413/5/ix1916/5 cmd[6] U9413/5/58 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-50.41 11.49 -50.28 11.64)
MU9413/5/ix1916/5 G_DG U9413/5/ix1916/SEL U9413/5/ix1916/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-49.83 11.49 -49.7 11.64)
MU9413/5/ix1916/6 U9413/5/ix1916/OUT U9413/5/58 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-49.25 11.49 -49.12 11.64)
MU9413/5/reg_r_shiftReg_51_/1 G_DG U9413/5/CLK U9413/5/42 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-66.475 11.49 -66.345 11.64)
MU9413/5/reg_r_shiftReg_51_/2 U9413/5/43 U9413/5/42 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-65.895 11.49 -65.765 11.64)
MU9413/5/reg_r_shiftReg_51_/3 U9413/5/reg_r_shiftReg_51_/4 U9413/5/ix1886/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-64.805 11.49 -64.675 11.64)
MU9413/5/reg_r_shiftReg_51_/4 U9413/5/46 U9413/5/42 U9413/5/reg_r_shiftReg_51_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-64.29 11.49 -64.16 11.64)
MU9413/5/reg_r_shiftReg_51_/5 U9413/5/47 U9413/5/46 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-63.2 11.49 -63.07 11.64)
MU9413/5/reg_r_shiftReg_51_/6 U9413/5/reg_r_shiftReg_51_/7 U9413/5/CLB U9413/5/46 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-61.83 11.49 -61.7 11.64)
MU9413/5/reg_r_shiftReg_51_/7 U9413/5/reg_r_shiftReg_51_/8 U9413/5/47 U9413/5/reg_r_shiftReg_51_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-61.35 11.49 -61.22 11.64)
MU9413/5/reg_r_shiftReg_51_/8 G_DG U9413/5/43 U9413/5/reg_r_shiftReg_51_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-60.87 11.49 -60.74 11.64)
MU9413/5/reg_r_shiftReg_51_/9 U9413/5/reg_r_shiftReg_51_/9 U9413/5/47 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-59.78 11.49 -59.65 11.64)
MU9413/5/reg_r_shiftReg_51_/10 U9413/5/reg_r_shiftReg_51_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_51_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-59.27 11.49 -59.14 11.64)
MU9413/5/reg_r_shiftReg_51_/11 U9413/5/50 U9413/5/43 U9413/5/reg_r_shiftReg_51_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-58.85 11.49 -58.72 11.64)
MU9413/5/reg_r_shiftReg_51_/12 U9413/5/51 U9413/5/50 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-57.76 11.49 -57.63 11.64)
MU9413/5/reg_r_shiftReg_51_/13 U9413/5/52 U9413/5/42 U9413/5/50 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-56.4 11.49 -56.27 11.64)
MU9413/5/reg_r_shiftReg_51_/14 U9413/5/reg_r_shiftReg_51_/14 U9413/5/CLB U9413/5/52 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-55.82 11.49 -55.69 11.64)
MU9413/5/reg_r_shiftReg_51_/15 G_DG U9413/5/51 U9413/5/reg_r_shiftReg_51_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-55.51 11.49 -55.38 11.64)
MU9413/5/reg_r_shiftReg_51_/16 cmd[6] U9413/5/52 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-54.42 11.49 -54.29 11.64)
MU9413/5/reg_r_shiftReg_51_/17 U9413/5/reg_r_shiftReg_51_/QB U9413/5/51 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-53.33 11.49 -53.2 11.64)
MU9413/5/ix1886/1 G_DG U9413/5/ix1876/SEL U9413/5/35 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-70.555 11.49 -70.425 11.64)
MU9413/5/ix1886/2 U9413/5/ix1886/3 U9413/5/35 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-69.975 11.49 -69.845 11.64)
MU9413/5/ix1886/3 U9413/5/37 cmd[6] U9413/5/ix1886/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-69.395 11.49 -69.265 11.64)
MU9413/5/ix1886/4 U9413/5/ix1886/5 cmd[5] U9413/5/37 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-68.815 11.49 -68.685 11.64)
MU9413/5/ix1886/5 G_DG U9413/5/ix1876/SEL U9413/5/ix1886/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-68.235 11.49 -68.105 11.64)
MU9413/5/ix1886/6 U9413/5/ix1886/OUT U9413/5/37 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-67.655 11.49 -67.525 11.64)
MU9413/5/reg_r_shiftReg_50_/1 G_DG U9413/5/CLK U9413/5/21 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-84.88 11.49 -84.75 11.64)
MU9413/5/reg_r_shiftReg_50_/2 U9413/5/22 U9413/5/21 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-84.3 11.49 -84.17 11.64)
MU9413/5/reg_r_shiftReg_50_/3 U9413/5/reg_r_shiftReg_50_/4 U9413/5/ix1876/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-83.21 11.49 -83.08 11.64)
MU9413/5/reg_r_shiftReg_50_/4 U9413/5/25 U9413/5/21 U9413/5/reg_r_shiftReg_50_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-82.695 11.49 -82.565 11.64)
MU9413/5/reg_r_shiftReg_50_/5 U9413/5/26 U9413/5/25 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-81.605 11.49 -81.475 11.64)
MU9413/5/reg_r_shiftReg_50_/6 U9413/5/reg_r_shiftReg_50_/7 U9413/5/CLB U9413/5/25 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-80.235 11.49 -80.105 11.64)
MU9413/5/reg_r_shiftReg_50_/7 U9413/5/reg_r_shiftReg_50_/8 U9413/5/26 U9413/5/reg_r_shiftReg_50_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-79.755 11.49 -79.625 11.64)
MU9413/5/reg_r_shiftReg_50_/8 G_DG U9413/5/22 U9413/5/reg_r_shiftReg_50_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-79.275 11.49 -79.145 11.64)
MU9413/5/reg_r_shiftReg_50_/9 U9413/5/reg_r_shiftReg_50_/9 U9413/5/26 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-78.185 11.49 -78.055 11.64)
MU9413/5/reg_r_shiftReg_50_/10 U9413/5/reg_r_shiftReg_50_/10 U9413/5/CLB U9413/5/reg_r_shiftReg_50_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-77.675 11.49 -77.545 11.64)
MU9413/5/reg_r_shiftReg_50_/11 U9413/5/29 U9413/5/22 U9413/5/reg_r_shiftReg_50_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-77.255 11.49 -77.125 11.64)
MU9413/5/reg_r_shiftReg_50_/12 U9413/5/30 U9413/5/29 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-76.165 11.49 -76.035 11.64)
MU9413/5/reg_r_shiftReg_50_/13 U9413/5/31 U9413/5/21 U9413/5/29 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-74.805 11.49 -74.675 11.64)
MU9413/5/reg_r_shiftReg_50_/14 U9413/5/reg_r_shiftReg_50_/14 U9413/5/CLB U9413/5/31 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-74.225 11.49 -74.095 11.64)
MU9413/5/reg_r_shiftReg_50_/15 G_DG U9413/5/30 U9413/5/reg_r_shiftReg_50_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-73.915 11.49 -73.785 11.64)
MU9413/5/reg_r_shiftReg_50_/16 cmd[5] U9413/5/31 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-72.825 11.49 -72.695 11.64)
MU9413/5/reg_r_shiftReg_50_/17 U9413/5/reg_r_shiftReg_50_/QB U9413/5/30 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-71.735 11.49 -71.605 11.64)
MU9413/5/ix1876/1 G_DG U9413/5/ix1876/SEL U9413/5/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-88.96 11.49 -88.83 11.64)
MU9413/5/ix1876/2 U9413/5/ix1876/3 U9413/5/14 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-88.38 11.49 -88.25 11.64)
MU9413/5/ix1876/3 U9413/5/16 cmd[5] U9413/5/ix1876/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-87.8 11.49 -87.67 11.64)
MU9413/5/ix1876/4 U9413/5/ix1876/5 cmd[4] U9413/5/16 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-87.22 11.49 -87.09 11.64)
MU9413/5/ix1876/5 G_DG U9413/5/ix1876/SEL U9413/5/ix1876/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-86.64 11.49 -86.51 11.64)
MU9413/5/ix1876/6 U9413/5/ix1876/OUT U9413/5/16 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-86.06 11.49 -85.93 11.64)
MU9413/5/ix1856/1 G_DG U9413/SEL U9413/5/6 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-93.04 11.49 -92.91 11.64)
MU9413/5/ix1856/2 U9413/5/ix1856/3 U9413/5/6 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-92.46 11.49 -92.33 11.64)
MU9413/5/ix1856/3 U9413/5/8 cmd[3] U9413/5/ix1856/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-91.88 11.49 -91.75 11.64)
MU9413/5/ix1856/4 U9413/5/ix1856/5 cmd[2] U9413/5/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-91.3 11.49 -91.17 11.64)
MU9413/5/ix1856/5 G_DG U9413/SEL U9413/5/ix1856/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-90.72 11.49 -90.59 11.64)
MU9413/5/ix1856/6 U9413/5/ix1856/OUT U9413/5/8 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-90.14 11.49 -90.01 11.64)
MU9413/6/1 G_DS CLK U9413/6/2 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-98.32 4.215 -98.19 4.515)
MU9413/6/2 U9413/6/CLK U9413/6/2 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-97.74 4.215 -97.61 4.515)
MU9413/6/3 G_DS CLK U9413/6/3 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-96.56 4.215 -96.43 4.515)
MU9413/6/4 U9413/6/CLK U9413/6/3 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-95.98 4.215 -95.85 4.515)
MU9413/6/5 G_DS CLK U9413/6/4 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-94.8 4.215 -94.67 4.515)
MU9413/6/6 U9413/6/CLK U9413/6/4 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-94.22 4.215 -94.09 4.515)
MU9413/6/7 G_DS U9413/6/CLK U9413/6/5 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-93.04 4.215 -92.91 4.515)
MU9413/6/8 U9413/6/6 U9413/6/5 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-92.46 4.215 -92.33 4.515)
MU9413/6/9 U9413/6/7 U9413/5/ix1856/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-91.37 4.215 -91.24 4.605)
MU9413/6/10 U9413/6/9 U9413/6/6 U9413/6/7 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-90.855 4.215 -90.725 4.605)
MU9413/6/11 U9413/6/10 U9413/6/9 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-89.765 4.215 -89.635 4.515)
MU9413/6/12 U9413/6/11 U9413/6/5 U9413/6/9 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-88.675 4.215 -88.545 4.605)
MU9413/6/13 G_DS U9413/6/CLB U9413/6/11 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-88.055 4.215 -87.925 4.605)
MU9413/6/14 U9413/6/11 U9413/6/10 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-87.435 4.215 -87.305 4.605)
MU9413/6/15 U9413/6/12 U9413/6/10 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-86.345 4.215 -86.215 4.605)
MU9413/6/16 U9413/6/13 U9413/6/5 U9413/6/12 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-86.035 4.215 -85.905 4.605)
MU9413/6/17 U9413/6/14 U9413/6/13 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-84.325 4.215 -84.195 4.515)
MU9413/6/18 U9413/6/15 U9413/6/6 U9413/6/13 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-83.235 4.215 -83.105 4.605)
MU9413/6/19 G_DS U9413/6/CLB U9413/6/15 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-82.655 4.215 -82.525 4.605)
MU9413/6/20 U9413/6/15 U9413/6/14 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-82.075 4.215 -81.945 4.515)
MU9413/6/21 cmd[3] U9413/6/15 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-80.985 4.215 -80.855 4.515)
MU9413/6/22 U9413/6/reg_r_shiftReg_48_/QB U9413/6/14 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-79.895 4.215 -79.765 4.515)
MU9413/6/23 G_DS U9413/5/ix1876/SEL U9413/6/19 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-78.715 4 -78.585 4.3)
MU9413/6/24 U9413/6/20 U9413/6/19 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-78.135 4 -78.005 4.52)
MU9413/6/25 U9413/6/21 cmd[3] U9413/6/20 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-77.555 4 -77.425 4.52)
MU9413/6/26 U9413/6/23 cmd[4] U9413/6/21 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-76.975 4 -76.845 4.52)
MU9413/6/27 G_DS U9413/5/ix1876/SEL U9413/6/23 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-76.395 4 -76.265 4.52)
MU9413/6/28 U9413/6/ix1866/OUT U9413/6/21 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-75.815 4.215 -75.685 4.515)
MU9413/6/29 G_DS U9413/6/CLK U9413/6/26 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-74.635 4.215 -74.505 4.515)
MU9413/6/30 U9413/6/27 U9413/6/26 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-74.055 4.215 -73.925 4.515)
MU9413/6/31 U9413/6/28 U9413/6/ix1866/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-72.965 4.215 -72.835 4.605)
MU9413/6/32 U9413/6/30 U9413/6/27 U9413/6/28 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-72.45 4.215 -72.32 4.605)
MU9413/6/33 U9413/6/31 U9413/6/30 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-71.36 4.215 -71.23 4.515)
MU9413/6/34 U9413/6/32 U9413/6/26 U9413/6/30 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-70.27 4.215 -70.14 4.605)
MU9413/6/35 G_DS U9413/6/CLB U9413/6/32 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-69.65 4.215 -69.52 4.605)
MU9413/6/36 U9413/6/32 U9413/6/31 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-69.03 4.215 -68.9 4.605)
MU9413/6/37 U9413/6/33 U9413/6/31 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-67.94 4.215 -67.81 4.605)
MU9413/6/38 U9413/6/34 U9413/6/26 U9413/6/33 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-67.63 4.215 -67.5 4.605)
MU9413/6/39 U9413/6/35 U9413/6/34 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-65.92 4.215 -65.79 4.515)
MU9413/6/40 U9413/6/36 U9413/6/27 U9413/6/34 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-64.83 4.215 -64.7 4.605)
MU9413/6/41 G_DS U9413/6/CLB U9413/6/36 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-64.25 4.215 -64.12 4.605)
MU9413/6/42 U9413/6/36 U9413/6/35 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-63.67 4.215 -63.54 4.515)
MU9413/6/43 cmd[4] U9413/6/36 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-62.58 4.215 -62.45 4.515)
MU9413/6/44 U9413/6/reg_r_shiftReg_49_/QB U9413/6/35 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-61.49 4.215 -61.36 4.515)
MU9413/6/45 G_DS U9413/6/CLK U9413/6/39 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-60.31 4.215 -60.18 4.515)
MU9413/6/46 U9413/6/40 U9413/6/39 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-59.73 4.215 -59.6 4.515)
MU9413/6/47 U9413/6/41 U9413/5/ix1916/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-58.64 4.215 -58.51 4.605)
MU9413/6/48 U9413/6/43 U9413/6/40 U9413/6/41 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-58.125 4.215 -57.995 4.605)
MU9413/6/49 U9413/6/44 U9413/6/43 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-57.035 4.215 -56.905 4.515)
MU9413/6/50 U9413/6/45 U9413/6/39 U9413/6/43 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-55.945 4.215 -55.815 4.605)
MU9413/6/51 G_DS U9413/6/CLB U9413/6/45 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-55.325 4.215 -55.195 4.605)
MU9413/6/52 U9413/6/45 U9413/6/44 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-54.705 4.215 -54.575 4.605)
MU9413/6/53 U9413/6/46 U9413/6/44 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-53.615 4.215 -53.485 4.605)
MU9413/6/54 U9413/6/47 U9413/6/39 U9413/6/46 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-53.305 4.215 -53.175 4.605)
MU9413/6/55 U9413/6/48 U9413/6/47 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-51.595 4.215 -51.465 4.515)
MU9413/6/56 U9413/6/49 U9413/6/40 U9413/6/47 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-50.505 4.215 -50.375 4.605)
MU9413/6/57 G_DS U9413/6/CLB U9413/6/49 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-49.925 4.215 -49.795 4.605)
MU9413/6/58 U9413/6/49 U9413/6/48 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-49.345 4.215 -49.215 4.515)
MU9413/6/59 readL U9413/6/49 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-48.255 4.215 -48.125 4.515)
MU9413/6/60 U9413/6/reg_r_readL/QB U9413/6/48 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-47.165 4.215 -47.035 4.515)
MU9413/6/61 G_DS U9413/5/ix1876/SEL U9413/6/53 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-45.985 4 -45.855 4.3)
MU9413/6/62 U9413/6/54 U9413/6/53 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-45.405 4 -45.275 4.52)
MU9413/6/63 U9413/6/55 U9413/5/ix1896/B U9413/6/54 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-44.825 4 -44.695 4.52)
MU9413/6/64 U9413/6/57 U9413/6/ix1926/B U9413/6/55 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-44.245 4 -44.115 4.52)
MU9413/6/65 G_DS U9413/5/ix1876/SEL U9413/6/57 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-43.665 4 -43.535 4.52)
MU9413/6/66 U9413/6/ix1926/OUT U9413/6/55 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-43.085 4.215 -42.955 4.515)
MU9413/6/67 G_DS U9413/6/CLK U9413/6/60 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-41.905 4.215 -41.775 4.515)
MU9413/6/68 U9413/6/61 U9413/6/60 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-41.325 4.215 -41.195 4.515)
MU9413/6/69 U9413/6/62 U9413/6/ix1926/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-40.235 4.215 -40.105 4.605)
MU9413/6/70 U9413/6/64 U9413/6/61 U9413/6/62 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-39.72 4.215 -39.59 4.605)
MU9413/6/71 U9413/6/65 U9413/6/64 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-38.63 4.215 -38.5 4.515)
MU9413/6/72 U9413/6/66 U9413/6/60 U9413/6/64 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-37.54 4.215 -37.41 4.605)
MU9413/6/73 G_DS U9413/6/CLB U9413/6/66 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-36.92 4.215 -36.79 4.605)
MU9413/6/74 U9413/6/66 U9413/6/65 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-36.3 4.215 -36.17 4.605)
MU9413/6/75 U9413/6/67 U9413/6/65 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-35.21 4.215 -35.08 4.605)
MU9413/6/76 U9413/6/68 U9413/6/60 U9413/6/67 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-34.9 4.215 -34.77 4.605)
MU9413/6/77 U9413/6/69 U9413/6/68 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-33.19 4.215 -33.06 4.515)
MU9413/6/78 U9413/6/70 U9413/6/61 U9413/6/68 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-32.1 4.215 -31.97 4.605)
MU9413/6/79 G_DS U9413/6/CLB U9413/6/70 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-31.52 4.215 -31.39 4.605)
MU9413/6/80 U9413/6/70 U9413/6/69 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-30.94 4.215 -30.81 4.515)
MU9413/6/81 U9413/6/ix1926/B U9413/6/70 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-29.85 4.215 -29.72 4.515)
MU9413/6/82 U9413/6/reg_r_shiftReg_53_/QB U9413/6/69 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-28.76 4.215 -28.63 4.515)
MU9413/6/83 G_DS U9413/5/ix1876/SEL U9413/6/74 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-27.58 4 -27.45 4.3)
MU9413/6/84 U9413/6/75 U9413/6/74 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-27 4 -26.87 4.52)
MU9413/6/85 U9413/6/76 U9413/6/ix1926/B U9413/6/75 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-26.42 4 -26.29 4.52)
MU9413/6/86 U9413/6/78 saciRsp U9413/6/76 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-25.84 4 -25.71 4.52)
MU9413/6/87 G_DS U9413/5/ix1876/SEL U9413/6/78 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-25.26 4 -25.13 4.52)
MU9413/6/88 U9413/6/ix1936/OUT U9413/6/76 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-24.68 4.215 -24.55 4.515)
MU9413/6/89 G_DS U9413/6/CLK U9413/6/81 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-23.5 4.215 -23.37 4.515)
MU9413/6/90 U9413/6/82 U9413/6/81 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-22.92 4.215 -22.79 4.515)
MU9413/6/91 U9413/6/83 U9413/6/ix1936/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(-21.83 4.215 -21.7 4.605)
MU9413/6/92 U9413/6/85 U9413/6/82 U9413/6/83 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(-21.315 4.215 -21.185 4.605)
MU9413/6/93 U9413/6/86 U9413/6/85 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-20.225 4.215 -20.095 4.515)
MU9413/6/94 U9413/6/87 U9413/6/81 U9413/6/85 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(-19.135 4.215 -19.005 4.605)
MU9413/6/95 G_DS U9413/6/CLB U9413/6/87 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(-18.515 4.215 -18.385 4.605)
MU9413/6/96 U9413/6/87 U9413/6/86 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(-17.895 4.215 -17.765 4.605)
MU9413/6/97 U9413/6/88 U9413/6/86 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(-16.805 4.215 -16.675 4.605)
MU9413/6/98 U9413/6/89 U9413/6/81 U9413/6/88 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(-16.495 4.215 -16.365 4.605)
MU9413/6/99 U9413/6/90 U9413/6/89 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-14.785 4.215 -14.655 4.515)
MU9413/6/100 U9413/6/91 U9413/6/82 U9413/6/89 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(-13.695 4.215 -13.565 4.605)
MU9413/6/101 G_DS U9413/6/CLB U9413/6/91 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(-13.115 4.215 -12.985 4.605)
MU9413/6/102 U9413/6/91 U9413/6/90 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(-12.535 4.215 -12.405 4.515)
MU9413/6/103 saciRsp U9413/6/91 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-11.445 4.215 -11.315 4.515)
MU9413/6/104 U9413/6/reg_r_shiftReg_54_/QB U9413/6/90 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(-10.355 4.215 -10.225 4.515)
MU9413/6/105 U9413/6/94 exec G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-9.175 4 -9.045 4.52)
MU9413/6/106 U9413/6/ix2000/OUT U9413/5/ix1896/B U9413/6/94 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-8.595 4 -8.465 4.52)
MU9413/6/107 U9413/6/98 ack G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=2.31e-013 ad=1.17e-013 pd=9.7e-007 ps=2.03e-006 nrd=0.432692 nrs=0.85429  $(-7.415 4 -7.285 4.52)
MU9413/6/108 U9413/6/ix1906/B U9413/6/ix2000/OUT U9413/6/98 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=2.31e-013 pd=2.03e-006 ps=9.7e-007 nrd=0.85429 nrs=0.432692  $(-6.835 4 -6.705 4.52)
MU9413/6/109 G_DS U9413/QB U9413/6/103 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(-5.655 4 -5.525 4.3)
MU9413/6/110 U9413/6/104 U9413/6/103 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(-5.075 4 -4.945 4.52)
MU9413/6/111 U9413/6/105 exec U9413/6/104 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(-4.495 4 -4.365 4.52)
MU9413/6/112 U9413/6/107 U9413/6/ix1906/B U9413/6/105 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(-3.915 4 -3.785 4.52)
MU9413/6/113 G_DS U9413/QB U9413/6/107 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(-3.335 4 -3.205 4.52)
MU9413/6/114 U9413/6/ix1906/OUT U9413/6/105 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(-2.755 4.215 -2.625 4.515)
MU9413/6/115 G_DS U9413/6/CLK U9413/6/110 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(-1.575 4.215 -1.445 4.515)
MU9413/6/116 U9413/6/111 U9413/6/110 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(-0.995 4.215 -0.865 4.515)
MU9413/6/117 U9413/6/112 U9413/6/ix1906/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(0.095 4.215 0.225 4.605)
MU9413/6/118 U9413/6/114 U9413/6/111 U9413/6/112 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(0.61 4.215 0.74 4.605)
MU9413/6/119 U9413/6/115 U9413/6/114 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(1.7 4.215 1.83 4.515)
MU9413/6/120 U9413/6/116 U9413/6/110 U9413/6/114 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(2.79 4.215 2.92 4.605)
MU9413/6/121 G_DS U9413/6/CLB U9413/6/116 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(3.41 4.215 3.54 4.605)
MU9413/6/122 U9413/6/116 U9413/6/115 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(4.03 4.215 4.16 4.605)
MU9413/6/123 U9413/6/117 U9413/6/115 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(5.12 4.215 5.25 4.605)
MU9413/6/124 U9413/6/118 U9413/6/110 U9413/6/117 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(5.43 4.215 5.56 4.605)
MU9413/6/125 U9413/6/119 U9413/6/118 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(7.14 4.215 7.27 4.515)
MU9413/6/126 U9413/6/120 U9413/6/111 U9413/6/118 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(8.23 4.215 8.36 4.605)
MU9413/6/127 G_DS U9413/6/CLB U9413/6/120 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(8.81 4.215 8.94 4.605)
MU9413/6/128 U9413/6/120 U9413/6/119 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(9.39 4.215 9.52 4.515)
MU9413/6/129 exec U9413/6/120 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(10.48 4.215 10.61 4.515)
MU9413/6/130 U9413/6/QB U9413/6/119 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(11.57 4.215 11.7 4.515)
MU9413/6/131 G_DS U9413/6/SEL U9413/6/123 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(12.75 4 12.88 4.3)
MU9413/6/132 U9413/6/124 U9413/6/123 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(13.33 4 13.46 4.52)
MU9413/6/133 U9413/6/125 U9413/6/ix1696/A U9413/6/124 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(13.91 4 14.04 4.52)
MU9413/6/134 U9413/6/127 U9413/4/ix2251/A U9413/6/125 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(14.49 4 14.62 4.52)
MU9413/6/135 G_DS U9413/6/SEL U9413/6/127 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(15.07 4 15.2 4.52)
MU9413/6/136 U9413/5/reg_r_shiftReg_0_/DATA U9413/6/125 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(15.65 4.215 15.78 4.515)
MU9413/6/137 U9413/6/ix2009/OUT U9413/6/CLK G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(16.83 4.215 16.96 4.515)
MU9413/6/138 G_DS U9413/6/ix2009/OUT U9413/6/132 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(18.01 4.215 18.14 4.515)
MU9413/6/139 U9413/6/133 U9413/6/132 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(18.59 4.215 18.72 4.515)
MU9413/6/140 U9413/6/134 saciCmd G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(19.68 4.215 19.81 4.605)
MU9413/6/141 U9413/6/136 U9413/6/133 U9413/6/134 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(20.195 4.215 20.325 4.605)
MU9413/6/142 U9413/6/137 U9413/6/136 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(21.285 4.215 21.415 4.515)
MU9413/6/143 U9413/6/138 U9413/6/132 U9413/6/136 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(22.375 4.215 22.505 4.605)
MU9413/6/144 G_DS U9413/6/CLB U9413/6/138 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(22.995 4.215 23.125 4.605)
MU9413/6/145 U9413/6/138 U9413/6/137 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(23.615 4.215 23.745 4.605)
MU9413/6/146 U9413/6/139 U9413/6/137 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(24.705 4.215 24.835 4.605)
MU9413/6/147 U9413/6/140 U9413/6/132 U9413/6/139 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(25.015 4.215 25.145 4.605)
MU9413/6/148 U9413/6/141 U9413/6/140 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(26.725 4.215 26.855 4.515)
MU9413/6/149 U9413/6/142 U9413/6/133 U9413/6/140 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(27.815 4.215 27.945 4.605)
MU9413/6/150 G_DS U9413/6/CLB U9413/6/142 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(28.395 4.215 28.525 4.605)
MU9413/6/151 U9413/6/142 U9413/6/141 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(28.975 4.215 29.105 4.515)
MU9413/6/152 U9413/6/ix1696/A U9413/6/142 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(30.065 4.215 30.195 4.515)
MU9413/6/153 U9413/6/reg_saciCmdFall/QB U9413/6/141 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(31.155 4.215 31.285 4.515)
MU9413/6/154 G_DS U9413/6/SEL U9413/6/146 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(32.335 4 32.465 4.3)
MU9413/6/155 U9413/6/147 U9413/6/146 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(32.915 4 33.045 4.52)
MU9413/6/156 U9413/6/148 wrData[31] U9413/6/147 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(33.495 4 33.625 4.52)
MU9413/6/157 U9413/6/150 addr[0] U9413/6/148 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(34.075 4 34.205 4.52)
MU9413/6/158 G_DS U9413/6/SEL U9413/6/150 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(34.655 4 34.785 4.52)
MU9413/6/159 U9413/6/ix1706/OUT U9413/6/148 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(35.235 4.215 35.365 4.515)
MU9413/6/160 G_DS U9413/6/CLK U9413/6/153 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(36.415 4.215 36.545 4.515)
MU9413/6/161 U9413/6/154 U9413/6/153 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(36.995 4.215 37.125 4.515)
MU9413/6/162 U9413/6/155 U9413/6/ix1706/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(38.085 4.215 38.215 4.605)
MU9413/6/163 U9413/6/157 U9413/6/154 U9413/6/155 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(38.6 4.215 38.73 4.605)
MU9413/6/164 U9413/6/158 U9413/6/157 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(39.69 4.215 39.82 4.515)
MU9413/6/165 U9413/6/159 U9413/6/153 U9413/6/157 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(40.78 4.215 40.91 4.605)
MU9413/6/166 G_DS U9413/6/CLB U9413/6/159 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(41.4 4.215 41.53 4.605)
MU9413/6/167 U9413/6/159 U9413/6/158 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(42.02 4.215 42.15 4.605)
MU9413/6/168 U9413/6/160 U9413/6/158 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(43.11 4.215 43.24 4.605)
MU9413/6/169 U9413/6/161 U9413/6/153 U9413/6/160 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(43.42 4.215 43.55 4.605)
MU9413/6/170 U9413/6/162 U9413/6/161 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(45.13 4.215 45.26 4.515)
MU9413/6/171 U9413/6/163 U9413/6/154 U9413/6/161 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(46.22 4.215 46.35 4.605)
MU9413/6/172 G_DS U9413/6/CLB U9413/6/163 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(46.8 4.215 46.93 4.605)
MU9413/6/173 U9413/6/163 U9413/6/162 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(47.38 4.215 47.51 4.515)
MU9413/6/174 addr[0] U9413/6/163 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(48.47 4.215 48.6 4.515)
MU9413/6/175 U9413/6/reg_r_shiftReg_33_/QB U9413/6/162 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(49.56 4.215 49.69 4.515)
MU9413/6/176 G_DS U9413/6/CLK U9413/6/166 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(50.74 4.215 50.87 4.515)
MU9413/6/177 U9413/6/167 U9413/6/166 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(51.32 4.215 51.45 4.515)
MU9413/6/178 U9413/6/168 U9413/5/ix1826/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(52.41 4.215 52.54 4.605)
MU9413/6/179 U9413/6/170 U9413/6/167 U9413/6/168 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(52.925 4.215 53.055 4.605)
MU9413/6/180 U9413/6/171 U9413/6/170 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(54.015 4.215 54.145 4.515)
MU9413/6/181 U9413/6/172 U9413/6/166 U9413/6/170 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(55.105 4.215 55.235 4.605)
MU9413/6/182 G_DS U9413/6/CLB U9413/6/172 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(55.725 4.215 55.855 4.605)
MU9413/6/183 U9413/6/172 U9413/6/171 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(56.345 4.215 56.475 4.605)
MU9413/6/184 U9413/6/173 U9413/6/171 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(57.435 4.215 57.565 4.605)
MU9413/6/185 U9413/6/174 U9413/6/166 U9413/6/173 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(57.745 4.215 57.875 4.605)
MU9413/6/186 U9413/6/175 U9413/6/174 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(59.455 4.215 59.585 4.515)
MU9413/6/187 U9413/6/176 U9413/6/167 U9413/6/174 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(60.545 4.215 60.675 4.605)
MU9413/6/188 G_DS U9413/6/CLB U9413/6/176 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(61.125 4.215 61.255 4.605)
MU9413/6/189 U9413/6/176 U9413/6/175 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(61.705 4.215 61.835 4.515)
MU9413/6/190 cmd[0] U9413/6/176 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(62.795 4.215 62.925 4.515)
MU9413/6/191 U9413/6/reg_r_shiftReg_45_/QB U9413/6/175 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(63.885 4.215 64.015 4.515)
MU9413/6/192 G_DS U9413/6/CLK U9413/6/179 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(65.065 4.215 65.195 4.515)
MU9413/6/193 U9413/6/180 U9413/6/179 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(65.645 4.215 65.775 4.515)
MU9413/6/194 U9413/6/181 U9413/reg_r_shiftReg_13_\Cross G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(66.735 4.215 66.865 4.605)
MU9413/6/195 U9413/6/183 U9413/6/180 U9413/6/181 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(67.25 4.215 67.38 4.605)
MU9413/6/196 U9413/6/184 U9413/6/183 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(68.34 4.215 68.47 4.515)
MU9413/6/197 U9413/6/185 U9413/6/179 U9413/6/183 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(69.43 4.215 69.56 4.605)
MU9413/6/198 G_DS U9413/6/CLB U9413/6/185 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(70.05 4.215 70.18 4.605)
MU9413/6/199 U9413/6/185 U9413/6/184 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(70.67 4.215 70.8 4.605)
MU9413/6/200 U9413/6/186 U9413/6/184 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(71.76 4.215 71.89 4.605)
MU9413/6/201 U9413/6/187 U9413/6/179 U9413/6/186 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(72.07 4.215 72.2 4.605)
MU9413/6/202 U9413/6/188 U9413/6/187 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(73.78 4.215 73.91 4.515)
MU9413/6/203 U9413/6/189 U9413/6/180 U9413/6/187 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(74.87 4.215 75 4.605)
MU9413/6/204 G_DS U9413/6/CLB U9413/6/189 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(75.45 4.215 75.58 4.605)
MU9413/6/205 U9413/6/189 U9413/6/188 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(76.03 4.215 76.16 4.515)
MU9413/6/206 wrData[8] U9413/6/189 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(77.12 4.215 77.25 4.515)
MU9413/6/207 U9413/6/reg_r_shiftReg_9_/QB U9413/6/188 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(78.21 4.215 78.34 4.515)
MU9413/6/208 G_DS U9413/6/SEL U9413/6/193 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(79.39 4 79.52 4.3)
MU9413/6/209 U9413/6/194 U9413/6/193 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(79.97 4 80.1 4.52)
MU9413/6/210 U9413/6/195 addr[0] U9413/6/194 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(80.55 4 80.68 4.52)
MU9413/6/211 U9413/6/197 addr[1] U9413/6/195 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(81.13 4 81.26 4.52)
MU9413/6/212 G_DS U9413/6/SEL U9413/6/197 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(81.71 4 81.84 4.52)
MU9413/6/213 U9413/6/ix1716/OUT U9413/6/195 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(82.29 4.215 82.42 4.515)
MU9413/6/214 G_DS U9413/6/SEL U9413/6/201 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(83.47 4 83.6 4.3)
MU9413/6/215 U9413/6/202 U9413/6/201 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(84.05 4 84.18 4.52)
MU9413/6/216 U9413/6/203 addr[1] U9413/6/202 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(84.63 4 84.76 4.52)
MU9413/6/217 U9413/6/205 addr[2] U9413/6/203 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(85.21 4 85.34 4.52)
MU9413/6/218 G_DS U9413/6/SEL U9413/6/205 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(85.79 4 85.92 4.52)
MU9413/6/219 U9413/5/reg_r_shiftReg_35_/DATA U9413/6/203 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(86.37 4.215 86.5 4.515)
MU9413/6/220 G_DS U9413/6/CLK U9413/6/208 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(87.55 4.215 87.68 4.515)
MU9413/6/221 U9413/6/209 U9413/6/208 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(88.13 4.215 88.26 4.515)
MU9413/6/222 U9413/6/210 U9413/6/ix1716/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(89.22 4.215 89.35 4.605)
MU9413/6/223 U9413/6/212 U9413/6/209 U9413/6/210 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(89.735 4.215 89.865 4.605)
MU9413/6/224 U9413/6/213 U9413/6/212 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(90.825 4.215 90.955 4.515)
MU9413/6/225 U9413/6/214 U9413/6/208 U9413/6/212 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(91.915 4.215 92.045 4.605)
MU9413/6/226 G_DS U9413/6/CLB U9413/6/214 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(92.535 4.215 92.665 4.605)
MU9413/6/227 U9413/6/214 U9413/6/213 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(93.155 4.215 93.285 4.605)
MU9413/6/228 U9413/6/215 U9413/6/213 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(94.245 4.215 94.375 4.605)
MU9413/6/229 U9413/6/216 U9413/6/208 U9413/6/215 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(94.555 4.215 94.685 4.605)
MU9413/6/230 U9413/6/217 U9413/6/216 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(96.265 4.215 96.395 4.515)
MU9413/6/231 U9413/6/218 U9413/6/209 U9413/6/216 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(97.355 4.215 97.485 4.605)
MU9413/6/232 G_DS U9413/6/CLB U9413/6/218 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(97.935 4.215 98.065 4.605)
MU9413/6/233 U9413/6/218 U9413/6/217 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(98.515 4.215 98.645 4.515)
MU9413/6/234 addr[1] U9413/6/218 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(99.605 4.215 99.735 4.515)
MU9413/6/235 U9413/6/reg_r_shiftReg_34_/QB U9413/6/217 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(100.695 4.215 100.825 4.515)
MU9413/6/236 G_DS U9413/6/SEL U9413/6/222 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(101.875 4 102.005 4.3)
MU9413/6/237 U9413/6/223 U9413/6/222 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(102.455 4 102.585 4.52)
MU9413/6/238 U9413/6/224 addr[2] U9413/6/223 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(103.035 4 103.165 4.52)
MU9413/6/239 U9413/6/226 addr[3] U9413/6/224 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(103.615 4 103.745 4.52)
MU9413/6/240 G_DS U9413/6/SEL U9413/6/226 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(104.195 4 104.325 4.52)
MU9413/6/241 U9413/6/ix1736/OUT U9413/6/224 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(104.775 4.215 104.905 4.515)
MU9413/6/242 G_DS U9413/6/CLK U9413/6/229 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(105.955 4.215 106.085 4.515)
MU9413/6/243 U9413/6/230 U9413/6/229 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(106.535 4.215 106.665 4.515)
MU9413/6/244 U9413/6/231 U9413/6/ix1736/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(107.625 4.215 107.755 4.605)
MU9413/6/245 U9413/6/233 U9413/6/230 U9413/6/231 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(108.14 4.215 108.27 4.605)
MU9413/6/246 U9413/6/234 U9413/6/233 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(109.23 4.215 109.36 4.515)
MU9413/6/247 U9413/6/235 U9413/6/229 U9413/6/233 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(110.32 4.215 110.45 4.605)
MU9413/6/248 G_DS U9413/6/CLB U9413/6/235 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(110.94 4.215 111.07 4.605)
MU9413/6/249 U9413/6/235 U9413/6/234 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(111.56 4.215 111.69 4.605)
MU9413/6/250 U9413/6/236 U9413/6/234 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(112.65 4.215 112.78 4.605)
MU9413/6/251 U9413/6/237 U9413/6/229 U9413/6/236 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(112.96 4.215 113.09 4.605)
MU9413/6/252 U9413/6/238 U9413/6/237 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(114.67 4.215 114.8 4.515)
MU9413/6/253 U9413/6/239 U9413/6/230 U9413/6/237 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(115.76 4.215 115.89 4.605)
MU9413/6/254 G_DS U9413/6/CLB U9413/6/239 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(116.34 4.215 116.47 4.605)
MU9413/6/255 U9413/6/239 U9413/6/238 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(116.92 4.215 117.05 4.515)
MU9413/6/256 addr[3] U9413/6/239 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(118.01 4.215 118.14 4.515)
MU9413/6/257 U9413/6/reg_r_shiftReg_36_/QB U9413/6/238 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(119.1 4.215 119.23 4.515)
MU9413/6/258 G_DS U9413/6/SEL U9413/6/243 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(120.28 4 120.41 4.3)
MU9413/6/259 U9413/6/244 U9413/6/243 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(120.86 4 120.99 4.52)
MU9413/6/260 U9413/6/245 addr[3] U9413/6/244 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(121.44 4 121.57 4.52)
MU9413/6/261 U9413/6/247 addr[4] U9413/6/245 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(122.02 4 122.15 4.52)
MU9413/6/262 G_DS U9413/6/SEL U9413/6/247 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(122.6 4 122.73 4.52)
MU9413/6/263 U9413/6/ix1746/OUT U9413/6/245 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(123.18 4.215 123.31 4.515)
MU9413/6/264 G_DS U9413/6/CLK U9413/6/250 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(124.36 4.215 124.49 4.515)
MU9413/6/265 U9413/6/251 U9413/6/250 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(124.94 4.215 125.07 4.515)
MU9413/6/266 U9413/6/252 U9413/6/ix1746/OUT G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(126.03 4.215 126.16 4.605)
MU9413/6/267 U9413/6/254 U9413/6/251 U9413/6/252 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(126.545 4.215 126.675 4.605)
MU9413/6/268 U9413/6/255 U9413/6/254 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(127.635 4.215 127.765 4.515)
MU9413/6/269 U9413/6/256 U9413/6/250 U9413/6/254 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(128.725 4.215 128.855 4.605)
MU9413/6/270 G_DS U9413/6/CLB U9413/6/256 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(129.345 4.215 129.475 4.605)
MU9413/6/271 U9413/6/256 U9413/6/255 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(129.965 4.215 130.095 4.605)
MU9413/6/272 U9413/6/257 U9413/6/255 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(131.055 4.215 131.185 4.605)
MU9413/6/273 U9413/6/258 U9413/6/250 U9413/6/257 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(131.365 4.215 131.495 4.605)
MU9413/6/274 U9413/6/259 U9413/6/258 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(133.075 4.215 133.205 4.515)
MU9413/6/275 U9413/6/260 U9413/6/251 U9413/6/258 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(134.165 4.215 134.295 4.605)
MU9413/6/276 G_DS U9413/6/CLB U9413/6/260 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(134.745 4.215 134.875 4.605)
MU9413/6/277 U9413/6/260 U9413/6/259 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(135.325 4.215 135.455 4.515)
MU9413/6/278 addr[4] U9413/6/260 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(136.415 4.215 136.545 4.515)
MU9413/6/279 U9413/6/reg_r_shiftReg_37_/QB U9413/6/259 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(137.505 4.215 137.635 4.515)
MU9413/6/280 G_DS U9413/6/SEL U9413/6/263 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=2.145e-013 ad=9.27439e-014 pd=7.97561e-007 ps=2.03e-006 nrd=1.03049 nrs=2.38333  $(138.685 4 138.815 4.3)
MU9413/6/281 U9413/6/264 U9413/6/263 G_DS G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.60756e-013 ad=1.17e-013 pd=9.7e-007 ps=1.38244e-006 nrd=0.432692 nrs=0.594512  $(139.265 4 139.395 4.52)
MU9413/6/282 U9413/6/265 addr[4] U9413/6/264 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.35e-013 pd=1.09e-006 ps=9.7e-007 nrd=0.49926 nrs=0.432692  $(139.845 4 139.975 4.52)
MU9413/6/283 U9413/6/266 addr[5] U9413/6/265 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.35e-013 ad=1.17e-013 pd=9.7e-007 ps=1.09e-006 nrd=0.432692 nrs=0.49926  $(140.425 4 140.555 4.52)
MU9413/6/284 G_DS U9413/6/SEL U9413/6/266 G_DS pch sa=-1 sb=-1 w=5.2e-007 l=1.3e-007 as=1.17e-013 ad=1.60756e-013 pd=1.38244e-006 ps=9.7e-007 nrd=0.594512 nrs=0.432692  $(141.005 4 141.135 4.52)
MU9413/6/285 U9413/6/DATA U9413/6/265 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=9.27439e-014 ad=1.395e-013 pd=1.53e-006 ps=7.97561e-007 nrd=1.55 nrs=1.03049  $(141.585 4.215 141.715 4.515)
MU9413/6/286 G_DS U9413/6/CLK U9413/6/267 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(142.765 4.215 142.895 4.515)
MU9413/6/287 U9413/6/268 U9413/6/267 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(143.345 4.215 143.475 4.515)
MU9413/6/288 U9413/6/269 U9413/6/DATA G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=7.5075e-014 pd=7.75e-007 ps=1.53e-006 nrd=0.49359 nrs=0.961538  $(144.435 4.215 144.565 4.605)
MU9413/6/289 U9413/6/270 U9413/6/268 U9413/6/269 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=7.5075e-014 ad=1.4625e-013 pd=1.53e-006 ps=7.75e-007 nrd=0.961538 nrs=0.49359  $(144.95 4.215 145.08 4.605)
MU9413/6/290 U9413/6/271 U9413/6/270 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(146.04 4.215 146.17 4.515)
MU9413/6/291 U9413/6/272 U9413/6/267 U9413/6/270 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=9.555e-014 pd=8.8e-007 ps=1.53e-006 nrd=0.628205 nrs=0.961538  $(147.13 4.215 147.26 4.605)
MU9413/6/292 G_DS U9413/6/CLB U9413/6/272 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=9.555e-014 pd=8.8e-007 ps=8.8e-007 nrd=0.628205 nrs=0.628205  $(147.75 4.215 147.88 4.605)
MU9413/6/293 U9413/6/272 U9413/6/271 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=9.555e-014 ad=1.4625e-013 pd=1.53e-006 ps=8.8e-007 nrd=0.961538 nrs=0.628205  $(148.37 4.215 148.5 4.605)
MU9413/6/294 U9413/6/273 U9413/6/271 G_DS G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=3.51e-014 pd=5.7e-007 ps=1.53e-006 nrd=0.230769 nrs=0.961538  $(149.46 4.215 149.59 4.605)
MU9413/6/295 U9413/6/274 U9413/6/267 U9413/6/273 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=3.51e-014 ad=1.4625e-013 pd=1.53e-006 ps=5.7e-007 nrd=0.961538 nrs=0.230769  $(149.77 4.215 149.9 4.605)
MU9413/6/296 U9413/6/275 U9413/6/274 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(151.48 4.215 151.61 4.515)
MU9413/6/297 U9413/6/276 U9413/6/268 U9413/6/274 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=1.4625e-013 ad=8.775e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.576923 nrs=0.961538  $(152.57 4.215 152.7 4.605)
MU9413/6/298 G_DS U9413/6/CLB U9413/6/276 G_DS pch sa=-1 sb=-1 w=3.9e-007 l=1.3e-007 as=8.775e-014 ad=9.53804e-014 pd=9.49565e-007 ps=8.4e-007 nrd=0.62709 nrs=0.576923  $(153.15 4.215 153.28 4.605)
MU9413/6/299 U9413/6/276 U9413/6/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=7.33696e-014 ad=1.395e-013 pd=1.53e-006 ps=7.30435e-007 nrd=1.55 nrs=0.815217  $(153.73 4.215 153.86 4.515)
MU9413/6/300 addr[5] U9413/6/276 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(154.82 4.215 154.95 4.515)
MU9413/6/301 U9413/6/reg_r_shiftReg_38_/QB U9413/6/275 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=1.395e-013 pd=1.53e-006 ps=1.53e-006 nrd=1.55 nrs=1.55  $(155.91 4.215 156.04 4.515)
MU9413/6/302 G_DS RST U9413/6/278 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(157.09 4.215 157.22 4.515)
MU9413/6/303 U9413/6/CLB U9413/6/278 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(157.67 4.215 157.8 4.515)
MU9413/6/304 G_DS RST U9413/6/279 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(158.85 4.215 158.98 4.515)
MU9413/6/305 U9413/6/CLB U9413/6/279 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(159.43 4.215 159.56 4.515)
MU9413/6/306 G_DS RST U9413/6/280 G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=1.395e-013 ad=8.1e-014 pd=8.4e-007 ps=1.53e-006 nrd=0.9 nrs=1.55  $(160.61 4.215 160.74 4.515)
MU9413/6/307 U9413/6/CLB U9413/6/280 G_DS G_DS pch sa=-1 sb=-1 w=3e-007 l=1.3e-007 as=8.1e-014 ad=1.395e-013 pd=1.53e-006 ps=8.4e-007 nrd=1.55 nrs=0.9  $(161.19 4.215 161.32 4.515)
MU9413/6/right_12/1 G_DG RST U9413/6/278 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(157.09 2.485 157.22 2.635)
MU9413/6/right_12/2 U9413/6/CLB U9413/6/278 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(157.67 2.485 157.8 2.635)
MU9413/6/right_11/1 G_DG RST U9413/6/279 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(158.85 2.485 158.98 2.635)
MU9413/6/right_11/2 U9413/6/CLB U9413/6/279 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(159.43 2.485 159.56 2.635)
MU9413/6/right_10/1 G_DG RST U9413/6/280 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(160.61 2.485 160.74 2.635)
MU9413/6/right_10/2 U9413/6/CLB U9413/6/280 G_DG G_DG nch sa=-2.15e-007 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(161.19 2.485 161.32 2.635)
MU9413/6/left_12/1 G_DG CLK U9413/6/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-96.56 2.485 -96.43 2.635)
MU9413/6/left_12/2 U9413/6/CLK U9413/6/3 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-95.98 2.485 -95.85 2.635)
MU9413/6/left_11/1 G_DG CLK U9413/6/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-94.8 2.485 -94.67 2.635)
MU9413/6/left_11/2 U9413/6/CLK U9413/6/4 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-94.22 2.485 -94.09 2.635)
MU9413/6/left_10/1 G_DG CLK U9413/6/2 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-98.32 2.485 -98.19 2.635)
MU9413/6/left_10/2 U9413/6/CLK U9413/6/2 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-97.74 2.485 -97.61 2.635)
MU9413/6/reg_r_shiftReg_38_/1 G_DG U9413/6/CLK U9413/6/267 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(142.765 2.485 142.895 2.635)
MU9413/6/reg_r_shiftReg_38_/2 U9413/6/268 U9413/6/267 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(143.345 2.485 143.475 2.635)
MU9413/6/reg_r_shiftReg_38_/3 U9413/6/reg_r_shiftReg_38_/4 U9413/6/DATA G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(144.435 2.485 144.565 2.635)
MU9413/6/reg_r_shiftReg_38_/4 U9413/6/270 U9413/6/267 U9413/6/reg_r_shiftReg_38_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(144.95 2.485 145.08 2.635)
MU9413/6/reg_r_shiftReg_38_/5 U9413/6/271 U9413/6/270 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(146.04 2.485 146.17 2.635)
MU9413/6/reg_r_shiftReg_38_/6 U9413/6/reg_r_shiftReg_38_/7 U9413/6/CLB U9413/6/270 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(147.41 2.485 147.54 2.635)
MU9413/6/reg_r_shiftReg_38_/7 U9413/6/reg_r_shiftReg_38_/8 U9413/6/271 U9413/6/reg_r_shiftReg_38_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(147.89 2.485 148.02 2.635)
MU9413/6/reg_r_shiftReg_38_/8 G_DG U9413/6/268 U9413/6/reg_r_shiftReg_38_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(148.37 2.485 148.5 2.635)
MU9413/6/reg_r_shiftReg_38_/9 U9413/6/reg_r_shiftReg_38_/9 U9413/6/271 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(149.46 2.485 149.59 2.635)
MU9413/6/reg_r_shiftReg_38_/10 U9413/6/reg_r_shiftReg_38_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_38_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(149.97 2.485 150.1 2.635)
MU9413/6/reg_r_shiftReg_38_/11 U9413/6/274 U9413/6/268 U9413/6/reg_r_shiftReg_38_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(150.39 2.485 150.52 2.635)
MU9413/6/reg_r_shiftReg_38_/12 U9413/6/275 U9413/6/274 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(151.48 2.485 151.61 2.635)
MU9413/6/reg_r_shiftReg_38_/13 U9413/6/276 U9413/6/267 U9413/6/274 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(152.84 2.485 152.97 2.635)
MU9413/6/reg_r_shiftReg_38_/14 U9413/6/reg_r_shiftReg_38_/14 U9413/6/CLB U9413/6/276 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(153.42 2.485 153.55 2.635)
MU9413/6/reg_r_shiftReg_38_/15 G_DG U9413/6/275 U9413/6/reg_r_shiftReg_38_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(153.73 2.485 153.86 2.635)
MU9413/6/reg_r_shiftReg_38_/16 addr[5] U9413/6/276 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(154.82 2.485 154.95 2.635)
MU9413/6/reg_r_shiftReg_38_/17 U9413/6/reg_r_shiftReg_38_/QB U9413/6/275 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(155.91 2.485 156.04 2.635)
MU9413/6/ix1756/1 G_DG U9413/6/SEL U9413/6/263 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(138.685 2.485 138.815 2.635)
MU9413/6/ix1756/2 U9413/6/ix1756/3 U9413/6/263 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(139.265 2.485 139.395 2.635)
MU9413/6/ix1756/3 U9413/6/265 addr[5] U9413/6/ix1756/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(139.845 2.485 139.975 2.635)
MU9413/6/ix1756/4 U9413/6/ix1756/5 addr[4] U9413/6/265 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(140.425 2.485 140.555 2.635)
MU9413/6/ix1756/5 G_DG U9413/6/SEL U9413/6/ix1756/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(141.005 2.485 141.135 2.635)
MU9413/6/ix1756/6 U9413/6/DATA U9413/6/265 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(141.585 2.485 141.715 2.635)
MU9413/6/reg_r_shiftReg_37_/1 G_DG U9413/6/CLK U9413/6/250 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(124.36 2.485 124.49 2.635)
MU9413/6/reg_r_shiftReg_37_/2 U9413/6/251 U9413/6/250 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(124.94 2.485 125.07 2.635)
MU9413/6/reg_r_shiftReg_37_/3 U9413/6/reg_r_shiftReg_37_/4 U9413/6/ix1746/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(126.03 2.485 126.16 2.635)
MU9413/6/reg_r_shiftReg_37_/4 U9413/6/254 U9413/6/250 U9413/6/reg_r_shiftReg_37_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(126.545 2.485 126.675 2.635)
MU9413/6/reg_r_shiftReg_37_/5 U9413/6/255 U9413/6/254 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(127.635 2.485 127.765 2.635)
MU9413/6/reg_r_shiftReg_37_/6 U9413/6/reg_r_shiftReg_37_/7 U9413/6/CLB U9413/6/254 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(129.005 2.485 129.135 2.635)
MU9413/6/reg_r_shiftReg_37_/7 U9413/6/reg_r_shiftReg_37_/8 U9413/6/255 U9413/6/reg_r_shiftReg_37_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(129.485 2.485 129.615 2.635)
MU9413/6/reg_r_shiftReg_37_/8 G_DG U9413/6/251 U9413/6/reg_r_shiftReg_37_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(129.965 2.485 130.095 2.635)
MU9413/6/reg_r_shiftReg_37_/9 U9413/6/reg_r_shiftReg_37_/9 U9413/6/255 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(131.055 2.485 131.185 2.635)
MU9413/6/reg_r_shiftReg_37_/10 U9413/6/reg_r_shiftReg_37_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_37_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(131.565 2.485 131.695 2.635)
MU9413/6/reg_r_shiftReg_37_/11 U9413/6/258 U9413/6/251 U9413/6/reg_r_shiftReg_37_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(131.985 2.485 132.115 2.635)
MU9413/6/reg_r_shiftReg_37_/12 U9413/6/259 U9413/6/258 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(133.075 2.485 133.205 2.635)
MU9413/6/reg_r_shiftReg_37_/13 U9413/6/260 U9413/6/250 U9413/6/258 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(134.435 2.485 134.565 2.635)
MU9413/6/reg_r_shiftReg_37_/14 U9413/6/reg_r_shiftReg_37_/14 U9413/6/CLB U9413/6/260 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(135.015 2.485 135.145 2.635)
MU9413/6/reg_r_shiftReg_37_/15 G_DG U9413/6/259 U9413/6/reg_r_shiftReg_37_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(135.325 2.485 135.455 2.635)
MU9413/6/reg_r_shiftReg_37_/16 addr[4] U9413/6/260 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(136.415 2.485 136.545 2.635)
MU9413/6/reg_r_shiftReg_37_/17 U9413/6/reg_r_shiftReg_37_/QB U9413/6/259 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(137.505 2.485 137.635 2.635)
MU9413/6/ix1746/1 G_DG U9413/6/SEL U9413/6/243 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(120.28 2.485 120.41 2.635)
MU9413/6/ix1746/2 U9413/6/ix1746/3 U9413/6/243 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(120.86 2.485 120.99 2.635)
MU9413/6/ix1746/3 U9413/6/245 addr[4] U9413/6/ix1746/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(121.44 2.485 121.57 2.635)
MU9413/6/ix1746/4 U9413/6/ix1746/5 addr[3] U9413/6/245 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(122.02 2.485 122.15 2.635)
MU9413/6/ix1746/5 G_DG U9413/6/SEL U9413/6/ix1746/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(122.6 2.485 122.73 2.635)
MU9413/6/ix1746/6 U9413/6/ix1746/OUT U9413/6/245 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(123.18 2.485 123.31 2.635)
MU9413/6/reg_r_shiftReg_36_/1 G_DG U9413/6/CLK U9413/6/229 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(105.955 2.485 106.085 2.635)
MU9413/6/reg_r_shiftReg_36_/2 U9413/6/230 U9413/6/229 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(106.535 2.485 106.665 2.635)
MU9413/6/reg_r_shiftReg_36_/3 U9413/6/reg_r_shiftReg_36_/4 U9413/6/ix1736/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(107.625 2.485 107.755 2.635)
MU9413/6/reg_r_shiftReg_36_/4 U9413/6/233 U9413/6/229 U9413/6/reg_r_shiftReg_36_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(108.14 2.485 108.27 2.635)
MU9413/6/reg_r_shiftReg_36_/5 U9413/6/234 U9413/6/233 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(109.23 2.485 109.36 2.635)
MU9413/6/reg_r_shiftReg_36_/6 U9413/6/reg_r_shiftReg_36_/7 U9413/6/CLB U9413/6/233 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(110.6 2.485 110.73 2.635)
MU9413/6/reg_r_shiftReg_36_/7 U9413/6/reg_r_shiftReg_36_/8 U9413/6/234 U9413/6/reg_r_shiftReg_36_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(111.08 2.485 111.21 2.635)
MU9413/6/reg_r_shiftReg_36_/8 G_DG U9413/6/230 U9413/6/reg_r_shiftReg_36_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(111.56 2.485 111.69 2.635)
MU9413/6/reg_r_shiftReg_36_/9 U9413/6/reg_r_shiftReg_36_/9 U9413/6/234 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(112.65 2.485 112.78 2.635)
MU9413/6/reg_r_shiftReg_36_/10 U9413/6/reg_r_shiftReg_36_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_36_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(113.16 2.485 113.29 2.635)
MU9413/6/reg_r_shiftReg_36_/11 U9413/6/237 U9413/6/230 U9413/6/reg_r_shiftReg_36_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(113.58 2.485 113.71 2.635)
MU9413/6/reg_r_shiftReg_36_/12 U9413/6/238 U9413/6/237 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(114.67 2.485 114.8 2.635)
MU9413/6/reg_r_shiftReg_36_/13 U9413/6/239 U9413/6/229 U9413/6/237 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(116.03 2.485 116.16 2.635)
MU9413/6/reg_r_shiftReg_36_/14 U9413/6/reg_r_shiftReg_36_/14 U9413/6/CLB U9413/6/239 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(116.61 2.485 116.74 2.635)
MU9413/6/reg_r_shiftReg_36_/15 G_DG U9413/6/238 U9413/6/reg_r_shiftReg_36_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(116.92 2.485 117.05 2.635)
MU9413/6/reg_r_shiftReg_36_/16 addr[3] U9413/6/239 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(118.01 2.485 118.14 2.635)
MU9413/6/reg_r_shiftReg_36_/17 U9413/6/reg_r_shiftReg_36_/QB U9413/6/238 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(119.1 2.485 119.23 2.635)
MU9413/6/ix1736/1 G_DG U9413/6/SEL U9413/6/222 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(101.875 2.485 102.005 2.635)
MU9413/6/ix1736/2 U9413/6/ix1736/3 U9413/6/222 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(102.455 2.485 102.585 2.635)
MU9413/6/ix1736/3 U9413/6/224 addr[3] U9413/6/ix1736/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(103.035 2.485 103.165 2.635)
MU9413/6/ix1736/4 U9413/6/ix1736/5 addr[2] U9413/6/224 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(103.615 2.485 103.745 2.635)
MU9413/6/ix1736/5 G_DG U9413/6/SEL U9413/6/ix1736/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(104.195 2.485 104.325 2.635)
MU9413/6/ix1736/6 U9413/6/ix1736/OUT U9413/6/224 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(104.775 2.485 104.905 2.635)
MU9413/6/reg_r_shiftReg_34_/1 G_DG U9413/6/CLK U9413/6/208 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(87.55 2.485 87.68 2.635)
MU9413/6/reg_r_shiftReg_34_/2 U9413/6/209 U9413/6/208 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(88.13 2.485 88.26 2.635)
MU9413/6/reg_r_shiftReg_34_/3 U9413/6/reg_r_shiftReg_34_/4 U9413/6/ix1716/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(89.22 2.485 89.35 2.635)
MU9413/6/reg_r_shiftReg_34_/4 U9413/6/212 U9413/6/208 U9413/6/reg_r_shiftReg_34_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(89.735 2.485 89.865 2.635)
MU9413/6/reg_r_shiftReg_34_/5 U9413/6/213 U9413/6/212 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(90.825 2.485 90.955 2.635)
MU9413/6/reg_r_shiftReg_34_/6 U9413/6/reg_r_shiftReg_34_/7 U9413/6/CLB U9413/6/212 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(92.195 2.485 92.325 2.635)
MU9413/6/reg_r_shiftReg_34_/7 U9413/6/reg_r_shiftReg_34_/8 U9413/6/213 U9413/6/reg_r_shiftReg_34_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(92.675 2.485 92.805 2.635)
MU9413/6/reg_r_shiftReg_34_/8 G_DG U9413/6/209 U9413/6/reg_r_shiftReg_34_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(93.155 2.485 93.285 2.635)
MU9413/6/reg_r_shiftReg_34_/9 U9413/6/reg_r_shiftReg_34_/9 U9413/6/213 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(94.245 2.485 94.375 2.635)
MU9413/6/reg_r_shiftReg_34_/10 U9413/6/reg_r_shiftReg_34_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_34_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(94.755 2.485 94.885 2.635)
MU9413/6/reg_r_shiftReg_34_/11 U9413/6/216 U9413/6/209 U9413/6/reg_r_shiftReg_34_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(95.175 2.485 95.305 2.635)
MU9413/6/reg_r_shiftReg_34_/12 U9413/6/217 U9413/6/216 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(96.265 2.485 96.395 2.635)
MU9413/6/reg_r_shiftReg_34_/13 U9413/6/218 U9413/6/208 U9413/6/216 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(97.625 2.485 97.755 2.635)
MU9413/6/reg_r_shiftReg_34_/14 U9413/6/reg_r_shiftReg_34_/14 U9413/6/CLB U9413/6/218 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(98.205 2.485 98.335 2.635)
MU9413/6/reg_r_shiftReg_34_/15 G_DG U9413/6/217 U9413/6/reg_r_shiftReg_34_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(98.515 2.485 98.645 2.635)
MU9413/6/reg_r_shiftReg_34_/16 addr[1] U9413/6/218 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(99.605 2.485 99.735 2.635)
MU9413/6/reg_r_shiftReg_34_/17 U9413/6/reg_r_shiftReg_34_/QB U9413/6/217 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(100.695 2.485 100.825 2.635)
MU9413/6/ix1726/1 G_DG U9413/6/SEL U9413/6/201 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(83.47 2.485 83.6 2.635)
MU9413/6/ix1726/2 U9413/6/ix1726/3 U9413/6/201 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(84.05 2.485 84.18 2.635)
MU9413/6/ix1726/3 U9413/6/203 addr[2] U9413/6/ix1726/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(84.63 2.485 84.76 2.635)
MU9413/6/ix1726/4 U9413/6/ix1726/5 addr[1] U9413/6/203 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(85.21 2.485 85.34 2.635)
MU9413/6/ix1726/5 G_DG U9413/6/SEL U9413/6/ix1726/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(85.79 2.485 85.92 2.635)
MU9413/6/ix1726/6 U9413/5/reg_r_shiftReg_35_/DATA U9413/6/203 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(86.37 2.485 86.5 2.635)
MU9413/6/ix1716/1 G_DG U9413/6/SEL U9413/6/193 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(79.39 2.485 79.52 2.635)
MU9413/6/ix1716/2 U9413/6/ix1716/3 U9413/6/193 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(79.97 2.485 80.1 2.635)
MU9413/6/ix1716/3 U9413/6/195 addr[1] U9413/6/ix1716/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(80.55 2.485 80.68 2.635)
MU9413/6/ix1716/4 U9413/6/ix1716/5 addr[0] U9413/6/195 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(81.13 2.485 81.26 2.635)
MU9413/6/ix1716/5 G_DG U9413/6/SEL U9413/6/ix1716/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(81.71 2.485 81.84 2.635)
MU9413/6/ix1716/6 U9413/6/ix1716/OUT U9413/6/195 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(82.29 2.485 82.42 2.635)
MU9413/6/reg_r_shiftReg_9_/1 G_DG U9413/6/CLK U9413/6/179 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(65.065 2.485 65.195 2.635)
MU9413/6/reg_r_shiftReg_9_/2 U9413/6/180 U9413/6/179 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(65.645 2.485 65.775 2.635)
MU9413/6/reg_r_shiftReg_9_/3 U9413/6/reg_r_shiftReg_9_/4 U9413/reg_r_shiftReg_13_\Cross G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(66.735 2.485 66.865 2.635)
MU9413/6/reg_r_shiftReg_9_/4 U9413/6/183 U9413/6/179 U9413/6/reg_r_shiftReg_9_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(67.25 2.485 67.38 2.635)
MU9413/6/reg_r_shiftReg_9_/5 U9413/6/184 U9413/6/183 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(68.34 2.485 68.47 2.635)
MU9413/6/reg_r_shiftReg_9_/6 U9413/6/reg_r_shiftReg_9_/7 U9413/6/CLB U9413/6/183 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(69.71 2.485 69.84 2.635)
MU9413/6/reg_r_shiftReg_9_/7 U9413/6/reg_r_shiftReg_9_/8 U9413/6/184 U9413/6/reg_r_shiftReg_9_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(70.19 2.485 70.32 2.635)
MU9413/6/reg_r_shiftReg_9_/8 G_DG U9413/6/180 U9413/6/reg_r_shiftReg_9_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(70.67 2.485 70.8 2.635)
MU9413/6/reg_r_shiftReg_9_/9 U9413/6/reg_r_shiftReg_9_/9 U9413/6/184 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(71.76 2.485 71.89 2.635)
MU9413/6/reg_r_shiftReg_9_/10 U9413/6/reg_r_shiftReg_9_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_9_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(72.27 2.485 72.4 2.635)
MU9413/6/reg_r_shiftReg_9_/11 U9413/6/187 U9413/6/180 U9413/6/reg_r_shiftReg_9_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(72.69 2.485 72.82 2.635)
MU9413/6/reg_r_shiftReg_9_/12 U9413/6/188 U9413/6/187 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(73.78 2.485 73.91 2.635)
MU9413/6/reg_r_shiftReg_9_/13 U9413/6/189 U9413/6/179 U9413/6/187 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(75.14 2.485 75.27 2.635)
MU9413/6/reg_r_shiftReg_9_/14 U9413/6/reg_r_shiftReg_9_/14 U9413/6/CLB U9413/6/189 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(75.72 2.485 75.85 2.635)
MU9413/6/reg_r_shiftReg_9_/15 G_DG U9413/6/188 U9413/6/reg_r_shiftReg_9_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(76.03 2.485 76.16 2.635)
MU9413/6/reg_r_shiftReg_9_/16 wrData[8] U9413/6/189 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(77.12 2.485 77.25 2.635)
MU9413/6/reg_r_shiftReg_9_/17 U9413/6/reg_r_shiftReg_9_/QB U9413/6/188 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(78.21 2.485 78.34 2.635)
MU9413/6/reg_r_shiftReg_45_/1 G_DG U9413/6/CLK U9413/6/166 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(50.74 2.485 50.87 2.635)
MU9413/6/reg_r_shiftReg_45_/2 U9413/6/167 U9413/6/166 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(51.32 2.485 51.45 2.635)
MU9413/6/reg_r_shiftReg_45_/3 U9413/6/reg_r_shiftReg_45_/4 U9413/5/ix1826/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(52.41 2.485 52.54 2.635)
MU9413/6/reg_r_shiftReg_45_/4 U9413/6/170 U9413/6/166 U9413/6/reg_r_shiftReg_45_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(52.925 2.485 53.055 2.635)
MU9413/6/reg_r_shiftReg_45_/5 U9413/6/171 U9413/6/170 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(54.015 2.485 54.145 2.635)
MU9413/6/reg_r_shiftReg_45_/6 U9413/6/reg_r_shiftReg_45_/7 U9413/6/CLB U9413/6/170 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(55.385 2.485 55.515 2.635)
MU9413/6/reg_r_shiftReg_45_/7 U9413/6/reg_r_shiftReg_45_/8 U9413/6/171 U9413/6/reg_r_shiftReg_45_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(55.865 2.485 55.995 2.635)
MU9413/6/reg_r_shiftReg_45_/8 G_DG U9413/6/167 U9413/6/reg_r_shiftReg_45_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(56.345 2.485 56.475 2.635)
MU9413/6/reg_r_shiftReg_45_/9 U9413/6/reg_r_shiftReg_45_/9 U9413/6/171 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(57.435 2.485 57.565 2.635)
MU9413/6/reg_r_shiftReg_45_/10 U9413/6/reg_r_shiftReg_45_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_45_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(57.945 2.485 58.075 2.635)
MU9413/6/reg_r_shiftReg_45_/11 U9413/6/174 U9413/6/167 U9413/6/reg_r_shiftReg_45_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(58.365 2.485 58.495 2.635)
MU9413/6/reg_r_shiftReg_45_/12 U9413/6/175 U9413/6/174 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(59.455 2.485 59.585 2.635)
MU9413/6/reg_r_shiftReg_45_/13 U9413/6/176 U9413/6/166 U9413/6/174 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(60.815 2.485 60.945 2.635)
MU9413/6/reg_r_shiftReg_45_/14 U9413/6/reg_r_shiftReg_45_/14 U9413/6/CLB U9413/6/176 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(61.395 2.485 61.525 2.635)
MU9413/6/reg_r_shiftReg_45_/15 G_DG U9413/6/175 U9413/6/reg_r_shiftReg_45_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(61.705 2.485 61.835 2.635)
MU9413/6/reg_r_shiftReg_45_/16 cmd[0] U9413/6/176 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(62.795 2.485 62.925 2.635)
MU9413/6/reg_r_shiftReg_45_/17 U9413/6/reg_r_shiftReg_45_/QB U9413/6/175 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(63.885 2.485 64.015 2.635)
MU9413/6/reg_r_shiftReg_33_/1 G_DG U9413/6/CLK U9413/6/153 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(36.415 2.485 36.545 2.635)
MU9413/6/reg_r_shiftReg_33_/2 U9413/6/154 U9413/6/153 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(36.995 2.485 37.125 2.635)
MU9413/6/reg_r_shiftReg_33_/3 U9413/6/reg_r_shiftReg_33_/4 U9413/6/ix1706/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(38.085 2.485 38.215 2.635)
MU9413/6/reg_r_shiftReg_33_/4 U9413/6/157 U9413/6/153 U9413/6/reg_r_shiftReg_33_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(38.6 2.485 38.73 2.635)
MU9413/6/reg_r_shiftReg_33_/5 U9413/6/158 U9413/6/157 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(39.69 2.485 39.82 2.635)
MU9413/6/reg_r_shiftReg_33_/6 U9413/6/reg_r_shiftReg_33_/7 U9413/6/CLB U9413/6/157 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(41.06 2.485 41.19 2.635)
MU9413/6/reg_r_shiftReg_33_/7 U9413/6/reg_r_shiftReg_33_/8 U9413/6/158 U9413/6/reg_r_shiftReg_33_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(41.54 2.485 41.67 2.635)
MU9413/6/reg_r_shiftReg_33_/8 G_DG U9413/6/154 U9413/6/reg_r_shiftReg_33_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(42.02 2.485 42.15 2.635)
MU9413/6/reg_r_shiftReg_33_/9 U9413/6/reg_r_shiftReg_33_/9 U9413/6/158 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(43.11 2.485 43.24 2.635)
MU9413/6/reg_r_shiftReg_33_/10 U9413/6/reg_r_shiftReg_33_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_33_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(43.62 2.485 43.75 2.635)
MU9413/6/reg_r_shiftReg_33_/11 U9413/6/161 U9413/6/154 U9413/6/reg_r_shiftReg_33_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(44.04 2.485 44.17 2.635)
MU9413/6/reg_r_shiftReg_33_/12 U9413/6/162 U9413/6/161 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(45.13 2.485 45.26 2.635)
MU9413/6/reg_r_shiftReg_33_/13 U9413/6/163 U9413/6/153 U9413/6/161 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(46.49 2.485 46.62 2.635)
MU9413/6/reg_r_shiftReg_33_/14 U9413/6/reg_r_shiftReg_33_/14 U9413/6/CLB U9413/6/163 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(47.07 2.485 47.2 2.635)
MU9413/6/reg_r_shiftReg_33_/15 G_DG U9413/6/162 U9413/6/reg_r_shiftReg_33_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(47.38 2.485 47.51 2.635)
MU9413/6/reg_r_shiftReg_33_/16 addr[0] U9413/6/163 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(48.47 2.485 48.6 2.635)
MU9413/6/reg_r_shiftReg_33_/17 U9413/6/reg_r_shiftReg_33_/QB U9413/6/162 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(49.56 2.485 49.69 2.635)
MU9413/6/ix1706/1 G_DG U9413/6/SEL U9413/6/146 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(32.335 2.485 32.465 2.635)
MU9413/6/ix1706/2 U9413/6/ix1706/3 U9413/6/146 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(32.915 2.485 33.045 2.635)
MU9413/6/ix1706/3 U9413/6/148 addr[0] U9413/6/ix1706/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(33.495 2.485 33.625 2.635)
MU9413/6/ix1706/4 U9413/6/ix1706/5 wrData[31] U9413/6/148 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(34.075 2.485 34.205 2.635)
MU9413/6/ix1706/5 G_DG U9413/6/SEL U9413/6/ix1706/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(34.655 2.485 34.785 2.635)
MU9413/6/ix1706/6 U9413/6/ix1706/OUT U9413/6/148 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(35.235 2.485 35.365 2.635)
MU9413/6/reg_saciCmdFall/1 G_DG U9413/6/ix2009/OUT U9413/6/132 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(18.01 2.485 18.14 2.635)
MU9413/6/reg_saciCmdFall/2 U9413/6/133 U9413/6/132 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(18.59 2.485 18.72 2.635)
MU9413/6/reg_saciCmdFall/3 U9413/6/reg_saciCmdFall/4 saciCmd G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(19.68 2.485 19.81 2.635)
MU9413/6/reg_saciCmdFall/4 U9413/6/136 U9413/6/132 U9413/6/reg_saciCmdFall/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(20.195 2.485 20.325 2.635)
MU9413/6/reg_saciCmdFall/5 U9413/6/137 U9413/6/136 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(21.285 2.485 21.415 2.635)
MU9413/6/reg_saciCmdFall/6 U9413/6/reg_saciCmdFall/7 U9413/6/CLB U9413/6/136 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(22.655 2.485 22.785 2.635)
MU9413/6/reg_saciCmdFall/7 U9413/6/reg_saciCmdFall/8 U9413/6/137 U9413/6/reg_saciCmdFall/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(23.135 2.485 23.265 2.635)
MU9413/6/reg_saciCmdFall/8 G_DG U9413/6/133 U9413/6/reg_saciCmdFall/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(23.615 2.485 23.745 2.635)
MU9413/6/reg_saciCmdFall/9 U9413/6/reg_saciCmdFall/9 U9413/6/137 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(24.705 2.485 24.835 2.635)
MU9413/6/reg_saciCmdFall/10 U9413/6/reg_saciCmdFall/10 U9413/6/CLB U9413/6/reg_saciCmdFall/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(25.215 2.485 25.345 2.635)
MU9413/6/reg_saciCmdFall/11 U9413/6/140 U9413/6/133 U9413/6/reg_saciCmdFall/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(25.635 2.485 25.765 2.635)
MU9413/6/reg_saciCmdFall/12 U9413/6/141 U9413/6/140 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(26.725 2.485 26.855 2.635)
MU9413/6/reg_saciCmdFall/13 U9413/6/142 U9413/6/132 U9413/6/140 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(28.085 2.485 28.215 2.635)
MU9413/6/reg_saciCmdFall/14 U9413/6/reg_saciCmdFall/14 U9413/6/CLB U9413/6/142 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(28.665 2.485 28.795 2.635)
MU9413/6/reg_saciCmdFall/15 G_DG U9413/6/141 U9413/6/reg_saciCmdFall/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(28.975 2.485 29.105 2.635)
MU9413/6/reg_saciCmdFall/16 U9413/6/ix1696/A U9413/6/142 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(30.065 2.485 30.195 2.635)
MU9413/6/reg_saciCmdFall/17 U9413/6/reg_saciCmdFall/QB U9413/6/141 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(31.155 2.485 31.285 2.635)
MU9413/6/ix2009/1 U9413/6/ix2009/OUT U9413/6/CLK G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(16.83 2.485 16.96 2.635)
MU9413/6/ix1696/1 G_DG U9413/6/SEL U9413/6/123 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(12.75 2.485 12.88 2.635)
MU9413/6/ix1696/2 U9413/6/ix1696/3 U9413/6/123 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(13.33 2.485 13.46 2.635)
MU9413/6/ix1696/3 U9413/6/125 U9413/4/ix2251/A U9413/6/ix1696/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(13.91 2.485 14.04 2.635)
MU9413/6/ix1696/4 U9413/6/ix1696/5 U9413/6/ix1696/A U9413/6/125 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(14.49 2.485 14.62 2.635)
MU9413/6/ix1696/5 G_DG U9413/6/SEL U9413/6/ix1696/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(15.07 2.485 15.2 2.635)
MU9413/6/ix1696/6 U9413/5/reg_r_shiftReg_0_/DATA U9413/6/125 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(15.65 2.485 15.78 2.635)
MU9413/6/reg_r_exec/1 G_DG U9413/6/CLK U9413/6/110 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-1.575 2.485 -1.445 2.635)
MU9413/6/reg_r_exec/2 U9413/6/111 U9413/6/110 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-0.995 2.485 -0.865 2.635)
MU9413/6/reg_r_exec/3 U9413/6/reg_r_exec/4 U9413/6/ix1906/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(0.095 2.485 0.225 2.635)
MU9413/6/reg_r_exec/4 U9413/6/114 U9413/6/110 U9413/6/reg_r_exec/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(0.61 2.485 0.74 2.635)
MU9413/6/reg_r_exec/5 U9413/6/115 U9413/6/114 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(1.7 2.485 1.83 2.635)
MU9413/6/reg_r_exec/6 U9413/6/reg_r_exec/7 U9413/6/CLB U9413/6/114 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(3.07 2.485 3.2 2.635)
MU9413/6/reg_r_exec/7 U9413/6/reg_r_exec/8 U9413/6/115 U9413/6/reg_r_exec/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(3.55 2.485 3.68 2.635)
MU9413/6/reg_r_exec/8 G_DG U9413/6/111 U9413/6/reg_r_exec/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(4.03 2.485 4.16 2.635)
MU9413/6/reg_r_exec/9 U9413/6/reg_r_exec/9 U9413/6/115 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(5.12 2.485 5.25 2.635)
MU9413/6/reg_r_exec/10 U9413/6/reg_r_exec/10 U9413/6/CLB U9413/6/reg_r_exec/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(5.63 2.485 5.76 2.635)
MU9413/6/reg_r_exec/11 U9413/6/118 U9413/6/111 U9413/6/reg_r_exec/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(6.05 2.485 6.18 2.635)
MU9413/6/reg_r_exec/12 U9413/6/119 U9413/6/118 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(7.14 2.485 7.27 2.635)
MU9413/6/reg_r_exec/13 U9413/6/120 U9413/6/110 U9413/6/118 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(8.5 2.485 8.63 2.635)
MU9413/6/reg_r_exec/14 U9413/6/reg_r_exec/14 U9413/6/CLB U9413/6/120 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(9.08 2.485 9.21 2.635)
MU9413/6/reg_r_exec/15 G_DG U9413/6/119 U9413/6/reg_r_exec/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(9.39 2.485 9.52 2.635)
MU9413/6/reg_r_exec/16 exec U9413/6/120 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(10.48 2.485 10.61 2.635)
MU9413/6/reg_r_exec/17 U9413/6/QB U9413/6/119 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(11.57 2.485 11.7 2.635)
MU9413/6/ix1906/1 G_DG U9413/QB U9413/6/103 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-5.655 2.485 -5.525 2.635)
MU9413/6/ix1906/2 U9413/6/ix1906/3 U9413/6/103 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-5.075 2.485 -4.945 2.635)
MU9413/6/ix1906/3 U9413/6/105 U9413/6/ix1906/B U9413/6/ix1906/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-4.495 2.485 -4.365 2.635)
MU9413/6/ix1906/4 U9413/6/ix1906/5 exec U9413/6/105 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-3.915 2.485 -3.785 2.635)
MU9413/6/ix1906/5 G_DG U9413/QB U9413/6/ix1906/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-3.335 2.485 -3.205 2.635)
MU9413/6/ix1906/6 U9413/6/ix1906/OUT U9413/6/105 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-2.755 2.485 -2.625 2.635)
MU9413/6/ix481/1 U9413/6/ix1906/B ack G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-7.415 2.485 -7.285 2.635)
MU9413/6/ix481/2 G_DG U9413/6/ix2000/OUT U9413/6/ix1906/B G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-6.835 2.485 -6.705 2.635)
MU9413/6/ix2000/1 U9413/6/ix2000/OUT exec G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-9.175 2.485 -9.045 2.635)
MU9413/6/ix2000/2 G_DG U9413/5/ix1896/B U9413/6/ix2000/OUT G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-8.595 2.485 -8.465 2.635)
MU9413/6/reg_r_shiftReg_54_/1 G_DG U9413/6/CLK U9413/6/81 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-23.5 2.485 -23.37 2.635)
MU9413/6/reg_r_shiftReg_54_/2 U9413/6/82 U9413/6/81 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-22.92 2.485 -22.79 2.635)
MU9413/6/reg_r_shiftReg_54_/3 U9413/6/reg_r_shiftReg_54_/4 U9413/6/ix1936/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-21.83 2.485 -21.7 2.635)
MU9413/6/reg_r_shiftReg_54_/4 U9413/6/85 U9413/6/81 U9413/6/reg_r_shiftReg_54_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-21.315 2.485 -21.185 2.635)
MU9413/6/reg_r_shiftReg_54_/5 U9413/6/86 U9413/6/85 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-20.225 2.485 -20.095 2.635)
MU9413/6/reg_r_shiftReg_54_/6 U9413/6/reg_r_shiftReg_54_/7 U9413/6/CLB U9413/6/85 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-18.855 2.485 -18.725 2.635)
MU9413/6/reg_r_shiftReg_54_/7 U9413/6/reg_r_shiftReg_54_/8 U9413/6/86 U9413/6/reg_r_shiftReg_54_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-18.375 2.485 -18.245 2.635)
MU9413/6/reg_r_shiftReg_54_/8 G_DG U9413/6/82 U9413/6/reg_r_shiftReg_54_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-17.895 2.485 -17.765 2.635)
MU9413/6/reg_r_shiftReg_54_/9 U9413/6/reg_r_shiftReg_54_/9 U9413/6/86 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-16.805 2.485 -16.675 2.635)
MU9413/6/reg_r_shiftReg_54_/10 U9413/6/reg_r_shiftReg_54_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_54_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-16.295 2.485 -16.165 2.635)
MU9413/6/reg_r_shiftReg_54_/11 U9413/6/89 U9413/6/82 U9413/6/reg_r_shiftReg_54_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-15.875 2.485 -15.745 2.635)
MU9413/6/reg_r_shiftReg_54_/12 U9413/6/90 U9413/6/89 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-14.785 2.485 -14.655 2.635)
MU9413/6/reg_r_shiftReg_54_/13 U9413/6/91 U9413/6/81 U9413/6/89 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-13.425 2.485 -13.295 2.635)
MU9413/6/reg_r_shiftReg_54_/14 U9413/6/reg_r_shiftReg_54_/14 U9413/6/CLB U9413/6/91 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-12.845 2.485 -12.715 2.635)
MU9413/6/reg_r_shiftReg_54_/15 G_DG U9413/6/90 U9413/6/reg_r_shiftReg_54_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-12.535 2.485 -12.405 2.635)
MU9413/6/reg_r_shiftReg_54_/16 saciRsp U9413/6/91 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-11.445 2.485 -11.315 2.635)
MU9413/6/reg_r_shiftReg_54_/17 U9413/6/reg_r_shiftReg_54_/QB U9413/6/90 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-10.355 2.485 -10.225 2.635)
MU9413/6/ix1936/1 G_DG U9413/5/ix1876/SEL U9413/6/74 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-27.58 2.485 -27.45 2.635)
MU9413/6/ix1936/2 U9413/6/ix1936/3 U9413/6/74 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-27 2.485 -26.87 2.635)
MU9413/6/ix1936/3 U9413/6/76 saciRsp U9413/6/ix1936/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-26.42 2.485 -26.29 2.635)
MU9413/6/ix1936/4 U9413/6/ix1936/5 U9413/6/ix1926/B U9413/6/76 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-25.84 2.485 -25.71 2.635)
MU9413/6/ix1936/5 G_DG U9413/5/ix1876/SEL U9413/6/ix1936/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-25.26 2.485 -25.13 2.635)
MU9413/6/ix1936/6 U9413/6/ix1936/OUT U9413/6/76 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-24.68 2.485 -24.55 2.635)
MU9413/6/reg_r_shiftReg_53_/1 G_DG U9413/6/CLK U9413/6/60 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-41.905 2.485 -41.775 2.635)
MU9413/6/reg_r_shiftReg_53_/2 U9413/6/61 U9413/6/60 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-41.325 2.485 -41.195 2.635)
MU9413/6/reg_r_shiftReg_53_/3 U9413/6/reg_r_shiftReg_53_/4 U9413/6/ix1926/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-40.235 2.485 -40.105 2.635)
MU9413/6/reg_r_shiftReg_53_/4 U9413/6/64 U9413/6/60 U9413/6/reg_r_shiftReg_53_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-39.72 2.485 -39.59 2.635)
MU9413/6/reg_r_shiftReg_53_/5 U9413/6/65 U9413/6/64 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-38.63 2.485 -38.5 2.635)
MU9413/6/reg_r_shiftReg_53_/6 U9413/6/reg_r_shiftReg_53_/7 U9413/6/CLB U9413/6/64 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-37.26 2.485 -37.13 2.635)
MU9413/6/reg_r_shiftReg_53_/7 U9413/6/reg_r_shiftReg_53_/8 U9413/6/65 U9413/6/reg_r_shiftReg_53_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-36.78 2.485 -36.65 2.635)
MU9413/6/reg_r_shiftReg_53_/8 G_DG U9413/6/61 U9413/6/reg_r_shiftReg_53_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-36.3 2.485 -36.17 2.635)
MU9413/6/reg_r_shiftReg_53_/9 U9413/6/reg_r_shiftReg_53_/9 U9413/6/65 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-35.21 2.485 -35.08 2.635)
MU9413/6/reg_r_shiftReg_53_/10 U9413/6/reg_r_shiftReg_53_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_53_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-34.7 2.485 -34.57 2.635)
MU9413/6/reg_r_shiftReg_53_/11 U9413/6/68 U9413/6/61 U9413/6/reg_r_shiftReg_53_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-34.28 2.485 -34.15 2.635)
MU9413/6/reg_r_shiftReg_53_/12 U9413/6/69 U9413/6/68 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-33.19 2.485 -33.06 2.635)
MU9413/6/reg_r_shiftReg_53_/13 U9413/6/70 U9413/6/60 U9413/6/68 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-31.83 2.485 -31.7 2.635)
MU9413/6/reg_r_shiftReg_53_/14 U9413/6/reg_r_shiftReg_53_/14 U9413/6/CLB U9413/6/70 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-31.25 2.485 -31.12 2.635)
MU9413/6/reg_r_shiftReg_53_/15 G_DG U9413/6/69 U9413/6/reg_r_shiftReg_53_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-30.94 2.485 -30.81 2.635)
MU9413/6/reg_r_shiftReg_53_/16 U9413/6/ix1926/B U9413/6/70 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-29.85 2.485 -29.72 2.635)
MU9413/6/reg_r_shiftReg_53_/17 U9413/6/reg_r_shiftReg_53_/QB U9413/6/69 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-28.76 2.485 -28.63 2.635)
MU9413/6/ix1926/1 G_DG U9413/5/ix1876/SEL U9413/6/53 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-45.985 2.485 -45.855 2.635)
MU9413/6/ix1926/2 U9413/6/ix1926/3 U9413/6/53 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-45.405 2.485 -45.275 2.635)
MU9413/6/ix1926/3 U9413/6/55 U9413/6/ix1926/B U9413/6/ix1926/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-44.825 2.485 -44.695 2.635)
MU9413/6/ix1926/4 U9413/6/ix1926/5 U9413/5/ix1896/B U9413/6/55 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-44.245 2.485 -44.115 2.635)
MU9413/6/ix1926/5 G_DG U9413/5/ix1876/SEL U9413/6/ix1926/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-43.665 2.485 -43.535 2.635)
MU9413/6/ix1926/6 U9413/6/ix1926/OUT U9413/6/55 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-43.085 2.485 -42.955 2.635)
MU9413/6/reg_r_readL/1 G_DG U9413/6/CLK U9413/6/39 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-60.31 2.485 -60.18 2.635)
MU9413/6/reg_r_readL/2 U9413/6/40 U9413/6/39 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-59.73 2.485 -59.6 2.635)
MU9413/6/reg_r_readL/3 U9413/6/reg_r_readL/4 U9413/5/ix1916/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-58.64 2.485 -58.51 2.635)
MU9413/6/reg_r_readL/4 U9413/6/43 U9413/6/39 U9413/6/reg_r_readL/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-58.125 2.485 -57.995 2.635)
MU9413/6/reg_r_readL/5 U9413/6/44 U9413/6/43 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-57.035 2.485 -56.905 2.635)
MU9413/6/reg_r_readL/6 U9413/6/reg_r_readL/7 U9413/6/CLB U9413/6/43 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-55.665 2.485 -55.535 2.635)
MU9413/6/reg_r_readL/7 U9413/6/reg_r_readL/8 U9413/6/44 U9413/6/reg_r_readL/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-55.185 2.485 -55.055 2.635)
MU9413/6/reg_r_readL/8 G_DG U9413/6/40 U9413/6/reg_r_readL/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-54.705 2.485 -54.575 2.635)
MU9413/6/reg_r_readL/9 U9413/6/reg_r_readL/9 U9413/6/44 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-53.615 2.485 -53.485 2.635)
MU9413/6/reg_r_readL/10 U9413/6/reg_r_readL/10 U9413/6/CLB U9413/6/reg_r_readL/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-53.105 2.485 -52.975 2.635)
MU9413/6/reg_r_readL/11 U9413/6/47 U9413/6/40 U9413/6/reg_r_readL/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-52.685 2.485 -52.555 2.635)
MU9413/6/reg_r_readL/12 U9413/6/48 U9413/6/47 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-51.595 2.485 -51.465 2.635)
MU9413/6/reg_r_readL/13 U9413/6/49 U9413/6/39 U9413/6/47 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-50.235 2.485 -50.105 2.635)
MU9413/6/reg_r_readL/14 U9413/6/reg_r_readL/14 U9413/6/CLB U9413/6/49 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-49.655 2.485 -49.525 2.635)
MU9413/6/reg_r_readL/15 G_DG U9413/6/48 U9413/6/reg_r_readL/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-49.345 2.485 -49.215 2.635)
MU9413/6/reg_r_readL/16 readL U9413/6/49 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-48.255 2.485 -48.125 2.635)
MU9413/6/reg_r_readL/17 U9413/6/reg_r_readL/QB U9413/6/48 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-47.165 2.485 -47.035 2.635)
MU9413/6/reg_r_shiftReg_49_/1 G_DG U9413/6/CLK U9413/6/26 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-74.635 2.485 -74.505 2.635)
MU9413/6/reg_r_shiftReg_49_/2 U9413/6/27 U9413/6/26 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-74.055 2.485 -73.925 2.635)
MU9413/6/reg_r_shiftReg_49_/3 U9413/6/reg_r_shiftReg_49_/4 U9413/6/ix1866/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-72.965 2.485 -72.835 2.635)
MU9413/6/reg_r_shiftReg_49_/4 U9413/6/30 U9413/6/26 U9413/6/reg_r_shiftReg_49_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-72.45 2.485 -72.32 2.635)
MU9413/6/reg_r_shiftReg_49_/5 U9413/6/31 U9413/6/30 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-71.36 2.485 -71.23 2.635)
MU9413/6/reg_r_shiftReg_49_/6 U9413/6/reg_r_shiftReg_49_/7 U9413/6/CLB U9413/6/30 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-69.99 2.485 -69.86 2.635)
MU9413/6/reg_r_shiftReg_49_/7 U9413/6/reg_r_shiftReg_49_/8 U9413/6/31 U9413/6/reg_r_shiftReg_49_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-69.51 2.485 -69.38 2.635)
MU9413/6/reg_r_shiftReg_49_/8 G_DG U9413/6/27 U9413/6/reg_r_shiftReg_49_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-69.03 2.485 -68.9 2.635)
MU9413/6/reg_r_shiftReg_49_/9 U9413/6/reg_r_shiftReg_49_/9 U9413/6/31 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-67.94 2.485 -67.81 2.635)
MU9413/6/reg_r_shiftReg_49_/10 U9413/6/reg_r_shiftReg_49_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_49_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-67.43 2.485 -67.3 2.635)
MU9413/6/reg_r_shiftReg_49_/11 U9413/6/34 U9413/6/27 U9413/6/reg_r_shiftReg_49_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-67.01 2.485 -66.88 2.635)
MU9413/6/reg_r_shiftReg_49_/12 U9413/6/35 U9413/6/34 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-65.92 2.485 -65.79 2.635)
MU9413/6/reg_r_shiftReg_49_/13 U9413/6/36 U9413/6/26 U9413/6/34 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-64.56 2.485 -64.43 2.635)
MU9413/6/reg_r_shiftReg_49_/14 U9413/6/reg_r_shiftReg_49_/14 U9413/6/CLB U9413/6/36 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-63.98 2.485 -63.85 2.635)
MU9413/6/reg_r_shiftReg_49_/15 G_DG U9413/6/35 U9413/6/reg_r_shiftReg_49_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-63.67 2.485 -63.54 2.635)
MU9413/6/reg_r_shiftReg_49_/16 cmd[4] U9413/6/36 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-62.58 2.485 -62.45 2.635)
MU9413/6/reg_r_shiftReg_49_/17 U9413/6/reg_r_shiftReg_49_/QB U9413/6/35 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-61.49 2.485 -61.36 2.635)
MU9413/6/ix1866/1 G_DG U9413/5/ix1876/SEL U9413/6/19 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-78.715 2.485 -78.585 2.635)
MU9413/6/ix1866/2 U9413/6/ix1866/3 U9413/6/19 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-78.135 2.485 -78.005 2.635)
MU9413/6/ix1866/3 U9413/6/21 cmd[4] U9413/6/ix1866/3 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-77.555 2.485 -77.425 2.635)
MU9413/6/ix1866/4 U9413/6/ix1866/5 cmd[3] U9413/6/21 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=3.375e-014 pd=6e-007 ps=8.6e-007 nrd=1.5 nrs=3.23333  $(-76.975 2.485 -76.845 2.635)
MU9413/6/ix1866/5 G_DG U9413/5/ix1876/SEL U9413/6/ix1866/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=3.375e-014 ad=7.275e-014 pd=8.6e-007 ps=6e-007 nrd=3.23333 nrs=1.5  $(-76.395 2.485 -76.265 2.635)
MU9413/6/ix1866/6 U9413/6/ix1866/OUT U9413/6/21 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-75.815 2.485 -75.685 2.635)
MU9413/6/reg_r_shiftReg_48_/1 G_DG U9413/6/CLK U9413/6/5 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-93.04 2.485 -92.91 2.635)
MU9413/6/reg_r_shiftReg_48_/2 U9413/6/6 U9413/6/5 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.3425e-013 pd=1.57e-006 ps=8.6e-007 nrd=5.96667 nrs=3.23333  $(-92.46 2.485 -92.33 2.635)
MU9413/6/reg_r_shiftReg_48_/3 U9413/6/reg_r_shiftReg_48_/4 U9413/5/ix1856/OUT G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.8875e-014 pd=5.35e-007 ps=1.57e-006 nrd=1.28333 nrs=5.96667  $(-91.37 2.485 -91.24 2.635)
MU9413/6/reg_r_shiftReg_48_/4 U9413/6/9 U9413/6/5 U9413/6/reg_r_shiftReg_48_/4 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.8875e-014 ad=1.3425e-013 pd=1.57e-006 ps=5.35e-007 nrd=5.96667 nrs=1.28333  $(-90.855 2.485 -90.725 2.635)
MU9413/6/reg_r_shiftReg_48_/5 U9413/6/10 U9413/6/9 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-89.765 2.485 -89.635 2.635)
MU9413/6/reg_r_shiftReg_48_/6 U9413/6/reg_r_shiftReg_48_/7 U9413/6/CLB U9413/6/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.625e-014 pd=5e-007 ps=1.57e-006 nrd=1.16667 nrs=5.96667  $(-88.395 2.485 -88.265 2.635)
MU9413/6/reg_r_shiftReg_48_/7 U9413/6/reg_r_shiftReg_48_/8 U9413/6/10 U9413/6/reg_r_shiftReg_48_/7 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=2.625e-014 pd=5e-007 ps=5e-007 nrd=1.16667 nrs=1.16667  $(-87.915 2.485 -87.785 2.635)
MU9413/6/reg_r_shiftReg_48_/8 G_DG U9413/6/6 U9413/6/reg_r_shiftReg_48_/8 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.625e-014 ad=1.3425e-013 pd=1.57e-006 ps=5e-007 nrd=5.96667 nrs=1.16667  $(-87.435 2.485 -87.305 2.635)
MU9413/6/reg_r_shiftReg_48_/9 U9413/6/reg_r_shiftReg_48_/9 U9413/6/10 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=2.85e-014 pd=5.3e-007 ps=1.57e-006 nrd=1.26667 nrs=5.96667  $(-86.345 2.485 -86.215 2.635)
MU9413/6/reg_r_shiftReg_48_/10 U9413/6/reg_r_shiftReg_48_/10 U9413/6/CLB U9413/6/reg_r_shiftReg_48_/9 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.85e-014 ad=2.175e-014 pd=4.4e-007 ps=5.3e-007 nrd=0.966667 nrs=1.26667  $(-85.835 2.485 -85.705 2.635)
MU9413/6/reg_r_shiftReg_48_/11 U9413/6/13 U9413/6/6 U9413/6/reg_r_shiftReg_48_/10 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=2.175e-014 ad=1.3425e-013 pd=1.57e-006 ps=4.4e-007 nrd=5.96667 nrs=0.966667  $(-85.415 2.485 -85.285 2.635)
MU9413/6/reg_r_shiftReg_48_/12 U9413/6/14 U9413/6/13 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-84.325 2.485 -84.195 2.635)
MU9413/6/reg_r_shiftReg_48_/13 U9413/6/15 U9413/6/5 U9413/6/13 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=7.275e-014 pd=8.6e-007 ps=1.57e-006 nrd=3.23333 nrs=5.96667  $(-82.965 2.485 -82.835 2.635)
MU9413/6/reg_r_shiftReg_48_/14 U9413/6/reg_r_shiftReg_48_/14 U9413/6/CLB U9413/6/15 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=7.275e-014 ad=1.35e-014 pd=3.3e-007 ps=8.6e-007 nrd=0.6 nrs=3.23333  $(-82.385 2.485 -82.255 2.635)
MU9413/6/reg_r_shiftReg_48_/15 G_DG U9413/6/14 U9413/6/reg_r_shiftReg_48_/14 G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.35e-014 ad=1.3425e-013 pd=1.57e-006 ps=3.3e-007 nrd=5.96667 nrs=0.6  $(-82.075 2.485 -81.945 2.635)
MU9413/6/reg_r_shiftReg_48_/16 cmd[3] U9413/6/15 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-80.985 2.485 -80.855 2.635)
MU9413/6/reg_r_shiftReg_48_/17 U9413/6/reg_r_shiftReg_48_/QB U9413/6/14 G_DG G_DG nch sa=-1 sb=-1 w=1.5e-007 l=1.3e-007 as=1.3425e-013 ad=1.3425e-013 pd=1.57e-006 ps=1.57e-006 nrd=5.96667 nrs=5.96667  $(-79.895 2.485 -79.765 2.635)

.ends
