../../saci/src/SaciSlaveWrapper.vhd