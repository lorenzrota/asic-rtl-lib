../../saci/src/saci_master.sv